* SPICE NETLIST
***************************************

.SUBCKT Eight_Bit_CSL_Adder VDD GND RESET CLK_MAIN SC0 SC1 SC2 SC3 SC4 SC5 SC6 SC7 C7_OUT S0 A0 B0 S1 A1 B1 S2
+ A2 B2 S3 A3 B3 S4 A4 B4 S5 A5 B5 S6 A6 B6 S7 A7 B7 Cout
** N=648 EP=38 IP=0 FDC=1276
M0 GND 5 S0 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.2e-14 AS=1.2e-14 PD=4.4e-07 PS=4.4e-07 $X=49850 $Y=49225 $D=1
M1 GND 10 248 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.2e-14 AS=1.2e-14 PD=4.4e-07 PS=4.4e-07 $X=50450 $Y=62980 $D=1
M2 GND 10 9 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.2e-14 AS=1.2e-14 PD=4.4e-07 PS=4.4e-07 $X=50450 $Y=63840 $D=1
M3 501 9 10 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.5e-14 AS=1.2e-14 PD=5e-07 PS=4.4e-07 $X=50450 $Y=64700 $D=1
M4 502 7 501 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.4e-14 AS=1.5e-14 PD=4.8e-07 PS=5e-07 $X=50450 $Y=65100 $D=1
M5 GND 4 502 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.2e-14 AS=1.4e-14 PD=4.4e-07 PS=4.8e-07 $X=50450 $Y=65480 $D=1
M6 GND RESET 7 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.2e-14 AS=1.2e-14 PD=4.4e-07 PS=4.4e-07 $X=50450 $Y=66360 $D=1
M7 GND 4 3 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.2e-14 AS=1.2e-14 PD=4.4e-07 PS=4.4e-07 $X=50450 $Y=67220 $D=1
M8 GND CLK_MAIN 4 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.2e-14 AS=1.2e-14 PD=4.4e-07 PS=4.4e-07 $X=50450 $Y=68080 $D=1
M9 11 3 10 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.2e-14 AS=1.2e-14 PD=4.4e-07 PS=4.4e-07 $X=50450 $Y=68940 $D=1
M10 503 3 GND GND NMOS_VTL L=5e-08 W=1e-07 AD=1.4e-14 AS=1.2e-14 PD=4.8e-07 PS=4.4e-07 $X=50450 $Y=69800 $D=1
M11 8 11 503 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.2e-14 AS=1.4e-14 PD=4.4e-07 PS=4.8e-07 $X=50450 $Y=70180 $D=1
M12 504 7 11 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.5e-14 AS=1.2e-14 PD=5e-07 PS=4.4e-07 $X=50450 $Y=71040 $D=1
M13 GND 8 504 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.2e-14 AS=1.5e-14 PD=4.4e-07 PS=5e-07 $X=50450 $Y=71440 $D=1
M14 249 4 8 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.2e-14 AS=1.2e-14 PD=4.4e-07 PS=4.4e-07 $X=50450 $Y=72300 $D=1
M15 GND 250 249 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.2e-14 AS=1.2e-14 PD=4.4e-07 PS=4.4e-07 $X=50450 $Y=73160 $D=1
M16 GND A0 250 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.2e-14 AS=1.2e-14 PD=4.4e-07 PS=4.4e-07 $X=50450 $Y=74020 $D=1
M17 GND 5 6 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.2e-14 AS=1.2e-14 PD=4.4e-07 PS=4.4e-07 $X=50710 $Y=49225 $D=1
M18 GND 248 252 GND NMOS_VTL L=5e-08 W=1.15e-07 AD=1.61e-14 AS=1.3225e-14 PD=5.1e-07 PS=4.6e-07 $X=50990 $Y=54715 $D=1
M19 GND 248 254 GND NMOS_VTL L=5e-08 W=1.15e-07 AD=1.61e-14 AS=1.3225e-14 PD=5.1e-07 PS=4.6e-07 $X=50990 $Y=57635 $D=1
M20 252 251 GND GND NMOS_VTL L=5e-08 W=1.15e-07 AD=1.61e-14 AS=1.61e-14 PD=5.1e-07 PS=5.1e-07 $X=51370 $Y=54715 $D=1
M21 254 251 GND GND NMOS_VTL L=5e-08 W=1.15e-07 AD=1.61e-14 AS=1.61e-14 PD=5.1e-07 PS=5.1e-07 $X=51370 $Y=57635 $D=1
M22 505 6 5 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.5e-14 AS=1.2e-14 PD=5e-07 PS=4.4e-07 $X=51570 $Y=49225 $D=1
M23 19 VDD 252 GND NMOS_VTL L=5e-08 W=1.15e-07 AD=1.61e-14 AS=1.61e-14 PD=5.1e-07 PS=5.1e-07 $X=51750 $Y=54715 $D=1
M24 20 GND 254 GND NMOS_VTL L=5e-08 W=1.15e-07 AD=1.61e-14 AS=1.61e-14 PD=5.1e-07 PS=5.1e-07 $X=51750 $Y=57635 $D=1
M25 506 17 505 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.4e-14 AS=1.5e-14 PD=4.8e-07 PS=5e-07 $X=51970 $Y=49225 $D=1
M26 507 248 19 GND NMOS_VTL L=5e-08 W=1.15e-07 AD=1.61e-14 AS=1.61e-14 PD=5.1e-07 PS=5.1e-07 $X=52130 $Y=54715 $D=1
M27 508 248 20 GND NMOS_VTL L=5e-08 W=1.15e-07 AD=1.61e-14 AS=1.61e-14 PD=5.1e-07 PS=5.1e-07 $X=52130 $Y=57635 $D=1
M28 GND 14 506 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.2e-14 AS=1.4e-14 PD=4.4e-07 PS=4.8e-07 $X=52350 $Y=49225 $D=1
M29 GND 251 507 GND NMOS_VTL L=5e-08 W=1.15e-07 AD=1.3225e-14 AS=1.61e-14 PD=4.6e-07 PS=5.1e-07 $X=52510 $Y=54715 $D=1
M30 GND 251 508 GND NMOS_VTL L=5e-08 W=1.15e-07 AD=1.3225e-14 AS=1.61e-14 PD=4.6e-07 PS=5.1e-07 $X=52510 $Y=57635 $D=1
M31 GND RESET 17 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.2e-14 AS=1.2e-14 PD=4.4e-07 PS=4.4e-07 $X=53230 $Y=49225 $D=1
M32 257 248 GND GND NMOS_VTL L=5e-08 W=1e-07 AD=1.4e-14 AS=1.15e-14 PD=4.8e-07 PS=4.3e-07 $X=53230 $Y=54745 $D=1
M33 259 248 GND GND NMOS_VTL L=5e-08 W=1e-07 AD=1.4e-14 AS=1.15e-14 PD=4.8e-07 PS=4.3e-07 $X=53230 $Y=57665 $D=1
M34 GND 251 257 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.4e-14 AS=1.4e-14 PD=4.8e-07 PS=4.8e-07 $X=53610 $Y=54745 $D=1
M35 GND 251 259 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.4e-14 AS=1.4e-14 PD=4.8e-07 PS=4.8e-07 $X=53610 $Y=57665 $D=1
M36 257 VDD GND GND NMOS_VTL L=5e-08 W=1e-07 AD=1.15e-14 AS=1.4e-14 PD=4.3e-07 PS=4.8e-07 $X=53990 $Y=54745 $D=1
M37 259 GND GND GND NMOS_VTL L=5e-08 W=1e-07 AD=1.15e-14 AS=1.4e-14 PD=4.3e-07 PS=4.8e-07 $X=53990 $Y=57665 $D=1
M38 GND 14 15 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.2e-14 AS=1.2e-14 PD=4.4e-07 PS=4.4e-07 $X=54090 $Y=49225 $D=1
M39 261 19 257 GND NMOS_VTL L=5e-08 W=9e-08 AD=1.08e-14 AS=1.125e-14 PD=4.2e-07 PS=4.3e-07 $X=54730 $Y=54745 $D=1
M40 262 20 259 GND NMOS_VTL L=5e-08 W=9e-08 AD=1.08e-14 AS=1.125e-14 PD=4.2e-07 PS=4.3e-07 $X=54730 $Y=57665 $D=1
M41 GND CLK_MAIN 14 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.2e-14 AS=1.2e-14 PD=4.4e-07 PS=4.4e-07 $X=54950 $Y=49225 $D=1
M42 509 VDD 261 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.4e-14 AS=1.15e-14 PD=4.8e-07 PS=4.3e-07 $X=55460 $Y=54745 $D=1
M43 510 GND 262 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.4e-14 AS=1.15e-14 PD=4.8e-07 PS=4.3e-07 $X=55460 $Y=57665 $D=1
M44 23 15 5 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.2e-14 AS=1.2e-14 PD=4.4e-07 PS=4.4e-07 $X=55810 $Y=49225 $D=1
M45 511 248 509 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.4e-14 AS=1.4e-14 PD=4.8e-07 PS=4.8e-07 $X=55840 $Y=54745 $D=1
M46 512 248 510 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.4e-14 AS=1.4e-14 PD=4.8e-07 PS=4.8e-07 $X=55840 $Y=57665 $D=1
M47 GND 27 251 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.2e-14 AS=1.2e-14 PD=4.4e-07 PS=4.4e-07 $X=55950 $Y=62980 $D=1
M48 GND 27 26 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.2e-14 AS=1.2e-14 PD=4.4e-07 PS=4.4e-07 $X=55950 $Y=63840 $D=1
M49 513 26 27 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.5e-14 AS=1.2e-14 PD=5e-07 PS=4.4e-07 $X=55950 $Y=64700 $D=1
M50 514 24 513 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.4e-14 AS=1.5e-14 PD=4.8e-07 PS=5e-07 $X=55950 $Y=65100 $D=1
M51 GND 22 514 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.2e-14 AS=1.4e-14 PD=4.4e-07 PS=4.8e-07 $X=55950 $Y=65480 $D=1
M52 GND RESET 24 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.2e-14 AS=1.2e-14 PD=4.4e-07 PS=4.4e-07 $X=55950 $Y=66360 $D=1
M53 GND 22 21 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.2e-14 AS=1.2e-14 PD=4.4e-07 PS=4.4e-07 $X=55950 $Y=67220 $D=1
M54 GND CLK_MAIN 22 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.2e-14 AS=1.2e-14 PD=4.4e-07 PS=4.4e-07 $X=55950 $Y=68080 $D=1
M55 28 21 27 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.2e-14 AS=1.2e-14 PD=4.4e-07 PS=4.4e-07 $X=55950 $Y=68940 $D=1
M56 515 21 GND GND NMOS_VTL L=5e-08 W=1e-07 AD=1.4e-14 AS=1.2e-14 PD=4.8e-07 PS=4.4e-07 $X=55950 $Y=69800 $D=1
M57 25 28 515 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.2e-14 AS=1.4e-14 PD=4.4e-07 PS=4.8e-07 $X=55950 $Y=70180 $D=1
M58 516 24 28 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.5e-14 AS=1.2e-14 PD=5e-07 PS=4.4e-07 $X=55950 $Y=71040 $D=1
M59 GND 25 516 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.2e-14 AS=1.5e-14 PD=4.4e-07 PS=5e-07 $X=55950 $Y=71440 $D=1
M60 263 22 25 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.2e-14 AS=1.2e-14 PD=4.4e-07 PS=4.4e-07 $X=55950 $Y=72300 $D=1
M61 GND 264 263 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.2e-14 AS=1.2e-14 PD=4.4e-07 PS=4.4e-07 $X=55950 $Y=73160 $D=1
M62 GND B0 264 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.2e-14 AS=1.2e-14 PD=4.4e-07 PS=4.4e-07 $X=55950 $Y=74020 $D=1
M63 GND 251 511 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.15e-14 AS=1.4e-14 PD=4.3e-07 PS=4.8e-07 $X=56220 $Y=54745 $D=1
M64 GND 251 512 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.15e-14 AS=1.4e-14 PD=4.3e-07 PS=4.8e-07 $X=56220 $Y=57665 $D=1
M65 517 15 GND GND NMOS_VTL L=5e-08 W=1e-07 AD=1.4e-14 AS=1.2e-14 PD=4.8e-07 PS=4.4e-07 $X=56670 $Y=49225 $D=1
M66 30 23 517 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.2e-14 AS=1.4e-14 PD=4.4e-07 PS=4.8e-07 $X=57050 $Y=49225 $D=1
M67 33 261 GND GND NMOS_VTL L=5e-08 W=1e-07 AD=1.2e-14 AS=1.2e-14 PD=4.4e-07 PS=4.4e-07 $X=57325 $Y=55295 $D=1
M68 266 GND GND GND NMOS_VTL L=5e-08 W=1e-07 AD=1.35e-14 AS=1.15e-14 PD=4.7e-07 PS=4.3e-07 $X=57350 $Y=57305 $D=1
M69 518 17 23 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.5e-14 AS=1.2e-14 PD=5e-07 PS=4.4e-07 $X=57910 $Y=49225 $D=1
M70 SC0 266 31 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.4e-14 AS=1.2e-14 PD=4.8e-07 PS=4.4e-07 $X=58120 $Y=57305 $D=1
M71 GND 30 518 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.2e-14 AS=1.5e-14 PD=4.4e-07 PS=5e-07 $X=58310 $Y=49225 $D=1
M72 GND 262 31 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.2e-14 AS=1.2e-14 PD=4.4e-07 PS=4.4e-07 $X=58330 $Y=58455 $D=1
M73 33 GND SC0 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.15e-14 AS=1.4e-14 PD=4.3e-07 PS=4.8e-07 $X=58500 $Y=57305 $D=1
M74 267 14 30 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.2e-14 AS=1.2e-14 PD=4.4e-07 PS=4.4e-07 $X=59170 $Y=49225 $D=1
M75 GND 268 267 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.2e-14 AS=1.2e-14 PD=4.4e-07 PS=4.4e-07 $X=60030 $Y=49225 $D=1
M76 GND SC0 268 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.2e-14 AS=1.2e-14 PD=4.4e-07 PS=4.4e-07 $X=60890 $Y=49225 $D=1
M77 GND 36 S1 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.2e-14 AS=1.2e-14 PD=4.4e-07 PS=4.4e-07 $X=62115 $Y=49225 $D=1
M78 GND 271 270 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.2e-14 AS=1.2e-14 PD=4.4e-07 PS=4.4e-07 $X=62155 $Y=61790 $D=1
M79 GND 41 271 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.2e-14 AS=1.2e-14 PD=4.4e-07 PS=4.4e-07 $X=62155 $Y=62975 $D=1
M80 GND 41 40 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.2e-14 AS=1.2e-14 PD=4.4e-07 PS=4.4e-07 $X=62155 $Y=63835 $D=1
M81 519 40 41 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.5e-14 AS=1.2e-14 PD=5e-07 PS=4.4e-07 $X=62155 $Y=64695 $D=1
M82 520 37 519 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.4e-14 AS=1.5e-14 PD=4.8e-07 PS=5e-07 $X=62155 $Y=65095 $D=1
M83 GND 35 520 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.2e-14 AS=1.4e-14 PD=4.4e-07 PS=4.8e-07 $X=62155 $Y=65475 $D=1
M84 GND RESET 37 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.2e-14 AS=1.2e-14 PD=4.4e-07 PS=4.4e-07 $X=62155 $Y=66355 $D=1
M85 GND 35 34 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.2e-14 AS=1.2e-14 PD=4.4e-07 PS=4.4e-07 $X=62155 $Y=67215 $D=1
M86 GND CLK_MAIN 35 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.2e-14 AS=1.2e-14 PD=4.4e-07 PS=4.4e-07 $X=62155 $Y=68075 $D=1
M87 42 34 41 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.2e-14 AS=1.2e-14 PD=4.4e-07 PS=4.4e-07 $X=62155 $Y=68935 $D=1
M88 521 34 GND GND NMOS_VTL L=5e-08 W=1e-07 AD=1.4e-14 AS=1.2e-14 PD=4.8e-07 PS=4.4e-07 $X=62155 $Y=69795 $D=1
M89 38 42 521 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.2e-14 AS=1.4e-14 PD=4.4e-07 PS=4.8e-07 $X=62155 $Y=70175 $D=1
M90 522 37 42 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.5e-14 AS=1.2e-14 PD=5e-07 PS=4.4e-07 $X=62155 $Y=71035 $D=1
M91 GND 38 522 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.2e-14 AS=1.5e-14 PD=4.4e-07 PS=5e-07 $X=62155 $Y=71435 $D=1
M92 272 35 38 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.2e-14 AS=1.2e-14 PD=4.4e-07 PS=4.4e-07 $X=62155 $Y=72295 $D=1
M93 GND 273 272 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.2e-14 AS=1.2e-14 PD=4.4e-07 PS=4.4e-07 $X=62155 $Y=73155 $D=1
M94 GND A1 273 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.2e-14 AS=1.2e-14 PD=4.4e-07 PS=4.4e-07 $X=62155 $Y=74015 $D=1
M95 GND 270 275 GND NMOS_VTL L=5e-08 W=1.15e-07 AD=1.61e-14 AS=1.3225e-14 PD=5.1e-07 PS=4.6e-07 $X=62790 $Y=54715 $D=1
M96 GND 270 277 GND NMOS_VTL L=5e-08 W=1.15e-07 AD=1.61e-14 AS=1.3225e-14 PD=5.1e-07 PS=4.6e-07 $X=62790 $Y=57795 $D=1
M97 GND 36 39 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.2e-14 AS=1.2e-14 PD=4.4e-07 PS=4.4e-07 $X=62975 $Y=49225 $D=1
M98 275 274 GND GND NMOS_VTL L=5e-08 W=1.15e-07 AD=1.61e-14 AS=1.61e-14 PD=5.1e-07 PS=5.1e-07 $X=63170 $Y=54715 $D=1
M99 277 274 GND GND NMOS_VTL L=5e-08 W=1.15e-07 AD=1.61e-14 AS=1.61e-14 PD=5.1e-07 PS=5.1e-07 $X=63170 $Y=57795 $D=1
M100 48 19 275 GND NMOS_VTL L=5e-08 W=1.15e-07 AD=1.61e-14 AS=1.61e-14 PD=5.1e-07 PS=5.1e-07 $X=63550 $Y=54715 $D=1
M101 49 20 277 GND NMOS_VTL L=5e-08 W=1.15e-07 AD=1.61e-14 AS=1.61e-14 PD=5.1e-07 PS=5.1e-07 $X=63550 $Y=57795 $D=1
M102 523 39 36 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.5e-14 AS=1.2e-14 PD=5e-07 PS=4.4e-07 $X=63835 $Y=49225 $D=1
M103 524 270 48 GND NMOS_VTL L=5e-08 W=1.15e-07 AD=1.61e-14 AS=1.61e-14 PD=5.1e-07 PS=5.1e-07 $X=63930 $Y=54715 $D=1
M104 525 270 49 GND NMOS_VTL L=5e-08 W=1.15e-07 AD=1.61e-14 AS=1.61e-14 PD=5.1e-07 PS=5.1e-07 $X=63930 $Y=57795 $D=1
M105 526 47 523 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.4e-14 AS=1.5e-14 PD=4.8e-07 PS=5e-07 $X=64235 $Y=49225 $D=1
M106 GND 274 524 GND NMOS_VTL L=5e-08 W=1.15e-07 AD=1.3225e-14 AS=1.61e-14 PD=4.6e-07 PS=5.1e-07 $X=64310 $Y=54715 $D=1
M107 GND 274 525 GND NMOS_VTL L=5e-08 W=1.15e-07 AD=1.3225e-14 AS=1.61e-14 PD=4.6e-07 PS=5.1e-07 $X=64310 $Y=57795 $D=1
M108 GND 45 526 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.2e-14 AS=1.4e-14 PD=4.4e-07 PS=4.8e-07 $X=64615 $Y=49225 $D=1
M109 280 270 GND GND NMOS_VTL L=5e-08 W=1e-07 AD=1.4e-14 AS=1.15e-14 PD=4.8e-07 PS=4.3e-07 $X=65030 $Y=54745 $D=1
M110 282 270 GND GND NMOS_VTL L=5e-08 W=1e-07 AD=1.4e-14 AS=1.15e-14 PD=4.8e-07 PS=4.3e-07 $X=65030 $Y=57825 $D=1
M111 GND 274 280 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.4e-14 AS=1.4e-14 PD=4.8e-07 PS=4.8e-07 $X=65410 $Y=54745 $D=1
M112 GND 274 282 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.4e-14 AS=1.4e-14 PD=4.8e-07 PS=4.8e-07 $X=65410 $Y=57825 $D=1
M113 GND RESET 47 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.2e-14 AS=1.2e-14 PD=4.4e-07 PS=4.4e-07 $X=65495 $Y=49225 $D=1
M114 280 19 GND GND NMOS_VTL L=5e-08 W=1e-07 AD=1.15e-14 AS=1.4e-14 PD=4.3e-07 PS=4.8e-07 $X=65790 $Y=54745 $D=1
M115 282 20 GND GND NMOS_VTL L=5e-08 W=1e-07 AD=1.15e-14 AS=1.4e-14 PD=4.3e-07 PS=4.8e-07 $X=65790 $Y=57825 $D=1
M116 GND 45 46 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.2e-14 AS=1.2e-14 PD=4.4e-07 PS=4.4e-07 $X=66355 $Y=49225 $D=1
M117 62 48 280 GND NMOS_VTL L=5e-08 W=9e-08 AD=1.08e-14 AS=1.125e-14 PD=4.2e-07 PS=4.3e-07 $X=66530 $Y=54745 $D=1
M118 60 49 282 GND NMOS_VTL L=5e-08 W=9e-08 AD=1.08e-14 AS=1.125e-14 PD=4.2e-07 PS=4.3e-07 $X=66530 $Y=57825 $D=1
M119 GND CLK_MAIN 45 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.2e-14 AS=1.2e-14 PD=4.4e-07 PS=4.4e-07 $X=67215 $Y=49225 $D=1
M120 527 19 62 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.4e-14 AS=1.15e-14 PD=4.8e-07 PS=4.3e-07 $X=67260 $Y=54745 $D=1
M121 528 20 60 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.4e-14 AS=1.15e-14 PD=4.8e-07 PS=4.3e-07 $X=67260 $Y=57825 $D=1
M122 533 270 527 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.4e-14 AS=1.4e-14 PD=4.8e-07 PS=4.8e-07 $X=67640 $Y=54745 $D=1
M123 534 270 528 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.4e-14 AS=1.4e-14 PD=4.8e-07 PS=4.8e-07 $X=67640 $Y=57825 $D=1
M124 GND 284 274 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.2e-14 AS=1.2e-14 PD=4.4e-07 PS=4.4e-07 $X=67675 $Y=61790 $D=1
M125 GND 55 284 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.2e-14 AS=1.2e-14 PD=4.4e-07 PS=4.4e-07 $X=67675 $Y=62975 $D=1
M126 GND 55 54 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.2e-14 AS=1.2e-14 PD=4.4e-07 PS=4.4e-07 $X=67675 $Y=63835 $D=1
M127 529 54 55 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.5e-14 AS=1.2e-14 PD=5e-07 PS=4.4e-07 $X=67675 $Y=64695 $D=1
M128 530 52 529 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.4e-14 AS=1.5e-14 PD=4.8e-07 PS=5e-07 $X=67675 $Y=65095 $D=1
M129 GND 51 530 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.2e-14 AS=1.4e-14 PD=4.4e-07 PS=4.8e-07 $X=67675 $Y=65475 $D=1
M130 GND RESET 52 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.2e-14 AS=1.2e-14 PD=4.4e-07 PS=4.4e-07 $X=67675 $Y=66355 $D=1
M131 GND 51 50 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.2e-14 AS=1.2e-14 PD=4.4e-07 PS=4.4e-07 $X=67675 $Y=67215 $D=1
M132 GND CLK_MAIN 51 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.2e-14 AS=1.2e-14 PD=4.4e-07 PS=4.4e-07 $X=67675 $Y=68075 $D=1
M133 56 50 55 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.2e-14 AS=1.2e-14 PD=4.4e-07 PS=4.4e-07 $X=67675 $Y=68935 $D=1
M134 531 50 GND GND NMOS_VTL L=5e-08 W=1e-07 AD=1.4e-14 AS=1.2e-14 PD=4.8e-07 PS=4.4e-07 $X=67675 $Y=69795 $D=1
M135 53 56 531 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.2e-14 AS=1.4e-14 PD=4.4e-07 PS=4.8e-07 $X=67675 $Y=70175 $D=1
M136 532 52 56 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.5e-14 AS=1.2e-14 PD=5e-07 PS=4.4e-07 $X=67675 $Y=71035 $D=1
M137 GND 53 532 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.2e-14 AS=1.5e-14 PD=4.4e-07 PS=5e-07 $X=67675 $Y=71435 $D=1
M138 285 51 53 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.2e-14 AS=1.2e-14 PD=4.4e-07 PS=4.4e-07 $X=67675 $Y=72295 $D=1
M139 GND 286 285 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.2e-14 AS=1.2e-14 PD=4.4e-07 PS=4.4e-07 $X=67675 $Y=73155 $D=1
M140 GND B1 286 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.2e-14 AS=1.2e-14 PD=4.4e-07 PS=4.4e-07 $X=67675 $Y=74015 $D=1
M141 GND 274 533 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.15e-14 AS=1.4e-14 PD=4.3e-07 PS=4.8e-07 $X=68020 $Y=54745 $D=1
M142 GND 274 534 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.15e-14 AS=1.4e-14 PD=4.3e-07 PS=4.8e-07 $X=68020 $Y=57825 $D=1
M143 57 46 36 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.2e-14 AS=1.2e-14 PD=4.4e-07 PS=4.4e-07 $X=68075 $Y=49225 $D=1
M144 535 46 GND GND NMOS_VTL L=5e-08 W=1e-07 AD=1.4e-14 AS=1.2e-14 PD=4.8e-07 PS=4.4e-07 $X=68935 $Y=49225 $D=1
M145 288 GND GND GND NMOS_VTL L=5e-08 W=1e-07 AD=1.35e-14 AS=1.15e-14 PD=4.7e-07 PS=4.3e-07 $X=69150 $Y=57465 $D=1
M146 59 57 535 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.2e-14 AS=1.4e-14 PD=4.4e-07 PS=4.8e-07 $X=69315 $Y=49225 $D=1
M147 SC1 288 60 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.4e-14 AS=1.2e-14 PD=4.8e-07 PS=4.4e-07 $X=69920 $Y=57465 $D=1
M148 536 47 57 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.5e-14 AS=1.2e-14 PD=5e-07 PS=4.4e-07 $X=70175 $Y=49225 $D=1
M149 62 GND SC1 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.15e-14 AS=1.4e-14 PD=4.3e-07 PS=4.8e-07 $X=70300 $Y=57465 $D=1
M150 GND 59 536 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.2e-14 AS=1.5e-14 PD=4.4e-07 PS=5e-07 $X=70575 $Y=49225 $D=1
M151 289 45 59 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.2e-14 AS=1.2e-14 PD=4.4e-07 PS=4.4e-07 $X=71435 $Y=49225 $D=1
M152 GND 290 289 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.2e-14 AS=1.2e-14 PD=4.4e-07 PS=4.4e-07 $X=72295 $Y=49225 $D=1
M153 GND SC1 290 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.2e-14 AS=1.2e-14 PD=4.4e-07 PS=4.4e-07 $X=73155 $Y=49225 $D=1
M154 GND 69 292 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.2e-14 AS=1.2e-14 PD=4.4e-07 PS=4.4e-07 $X=74050 $Y=62980 $D=1
M155 GND 69 68 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.2e-14 AS=1.2e-14 PD=4.4e-07 PS=4.4e-07 $X=74050 $Y=63840 $D=1
M156 537 68 69 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.5e-14 AS=1.2e-14 PD=5e-07 PS=4.4e-07 $X=74050 $Y=64700 $D=1
M157 538 65 537 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.4e-14 AS=1.5e-14 PD=4.8e-07 PS=5e-07 $X=74050 $Y=65100 $D=1
M158 GND 64 538 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.2e-14 AS=1.4e-14 PD=4.4e-07 PS=4.8e-07 $X=74050 $Y=65480 $D=1
M159 GND RESET 65 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.2e-14 AS=1.2e-14 PD=4.4e-07 PS=4.4e-07 $X=74050 $Y=66360 $D=1
M160 GND 64 63 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.2e-14 AS=1.2e-14 PD=4.4e-07 PS=4.4e-07 $X=74050 $Y=67220 $D=1
M161 GND CLK_MAIN 64 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.2e-14 AS=1.2e-14 PD=4.4e-07 PS=4.4e-07 $X=74050 $Y=68080 $D=1
M162 70 63 69 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.2e-14 AS=1.2e-14 PD=4.4e-07 PS=4.4e-07 $X=74050 $Y=68940 $D=1
M163 539 63 GND GND NMOS_VTL L=5e-08 W=1e-07 AD=1.4e-14 AS=1.2e-14 PD=4.8e-07 PS=4.4e-07 $X=74050 $Y=69800 $D=1
M164 66 70 539 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.2e-14 AS=1.4e-14 PD=4.4e-07 PS=4.8e-07 $X=74050 $Y=70180 $D=1
M165 540 65 70 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.5e-14 AS=1.2e-14 PD=5e-07 PS=4.4e-07 $X=74050 $Y=71040 $D=1
M166 GND 66 540 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.2e-14 AS=1.5e-14 PD=4.4e-07 PS=5e-07 $X=74050 $Y=71440 $D=1
M167 293 64 66 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.2e-14 AS=1.2e-14 PD=4.4e-07 PS=4.4e-07 $X=74050 $Y=72300 $D=1
M168 GND 294 293 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.2e-14 AS=1.2e-14 PD=4.4e-07 PS=4.4e-07 $X=74050 $Y=73160 $D=1
M169 GND A2 294 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.2e-14 AS=1.2e-14 PD=4.4e-07 PS=4.4e-07 $X=74050 $Y=74020 $D=1
M170 GND 67 S2 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.2e-14 AS=1.2e-14 PD=4.4e-07 PS=4.4e-07 $X=74310 $Y=49225 $D=1
M171 GND 292 296 GND NMOS_VTL L=5e-08 W=1.15e-07 AD=1.61e-14 AS=1.3225e-14 PD=5.1e-07 PS=4.6e-07 $X=74590 $Y=54715 $D=1
M172 GND 292 298 GND NMOS_VTL L=5e-08 W=1.15e-07 AD=1.61e-14 AS=1.3225e-14 PD=5.1e-07 PS=4.6e-07 $X=74590 $Y=57795 $D=1
M173 296 295 GND GND NMOS_VTL L=5e-08 W=1.15e-07 AD=1.61e-14 AS=1.61e-14 PD=5.1e-07 PS=5.1e-07 $X=74970 $Y=54715 $D=1
M174 298 295 GND GND NMOS_VTL L=5e-08 W=1.15e-07 AD=1.61e-14 AS=1.61e-14 PD=5.1e-07 PS=5.1e-07 $X=74970 $Y=57795 $D=1
M175 GND 67 71 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.2e-14 AS=1.2e-14 PD=4.4e-07 PS=4.4e-07 $X=75170 $Y=49225 $D=1
M176 77 48 296 GND NMOS_VTL L=5e-08 W=1.15e-07 AD=1.61e-14 AS=1.61e-14 PD=5.1e-07 PS=5.1e-07 $X=75350 $Y=54715 $D=1
M177 78 49 298 GND NMOS_VTL L=5e-08 W=1.15e-07 AD=1.61e-14 AS=1.61e-14 PD=5.1e-07 PS=5.1e-07 $X=75350 $Y=57795 $D=1
M178 541 292 77 GND NMOS_VTL L=5e-08 W=1.15e-07 AD=1.61e-14 AS=1.61e-14 PD=5.1e-07 PS=5.1e-07 $X=75730 $Y=54715 $D=1
M179 542 292 78 GND NMOS_VTL L=5e-08 W=1.15e-07 AD=1.61e-14 AS=1.61e-14 PD=5.1e-07 PS=5.1e-07 $X=75730 $Y=57795 $D=1
M180 543 71 67 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.5e-14 AS=1.2e-14 PD=5e-07 PS=4.4e-07 $X=76030 $Y=49225 $D=1
M181 GND 295 541 GND NMOS_VTL L=5e-08 W=1.15e-07 AD=1.3225e-14 AS=1.61e-14 PD=4.6e-07 PS=5.1e-07 $X=76110 $Y=54715 $D=1
M182 GND 295 542 GND NMOS_VTL L=5e-08 W=1.15e-07 AD=1.3225e-14 AS=1.61e-14 PD=4.6e-07 PS=5.1e-07 $X=76110 $Y=57795 $D=1
M183 544 76 543 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.4e-14 AS=1.5e-14 PD=4.8e-07 PS=5e-07 $X=76430 $Y=49225 $D=1
M184 GND 74 544 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.2e-14 AS=1.4e-14 PD=4.4e-07 PS=4.8e-07 $X=76810 $Y=49225 $D=1
M185 301 292 GND GND NMOS_VTL L=5e-08 W=1e-07 AD=1.4e-14 AS=1.15e-14 PD=4.8e-07 PS=4.3e-07 $X=76830 $Y=54745 $D=1
M186 303 292 GND GND NMOS_VTL L=5e-08 W=1e-07 AD=1.4e-14 AS=1.15e-14 PD=4.8e-07 PS=4.3e-07 $X=76830 $Y=57825 $D=1
M187 GND 295 301 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.4e-14 AS=1.4e-14 PD=4.8e-07 PS=4.8e-07 $X=77210 $Y=54745 $D=1
M188 GND 295 303 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.4e-14 AS=1.4e-14 PD=4.8e-07 PS=4.8e-07 $X=77210 $Y=57825 $D=1
M189 301 48 GND GND NMOS_VTL L=5e-08 W=1e-07 AD=1.15e-14 AS=1.4e-14 PD=4.3e-07 PS=4.8e-07 $X=77590 $Y=54745 $D=1
M190 303 49 GND GND NMOS_VTL L=5e-08 W=1e-07 AD=1.15e-14 AS=1.4e-14 PD=4.3e-07 PS=4.8e-07 $X=77590 $Y=57825 $D=1
M191 GND RESET 76 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.2e-14 AS=1.2e-14 PD=4.4e-07 PS=4.4e-07 $X=77690 $Y=49225 $D=1
M192 305 77 301 GND NMOS_VTL L=5e-08 W=9e-08 AD=1.08e-14 AS=1.125e-14 PD=4.2e-07 PS=4.3e-07 $X=78330 $Y=54745 $D=1
M193 306 78 303 GND NMOS_VTL L=5e-08 W=9e-08 AD=1.08e-14 AS=1.125e-14 PD=4.2e-07 PS=4.3e-07 $X=78330 $Y=57825 $D=1
M194 GND 74 75 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.2e-14 AS=1.2e-14 PD=4.4e-07 PS=4.4e-07 $X=78550 $Y=49225 $D=1
M195 545 48 305 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.4e-14 AS=1.15e-14 PD=4.8e-07 PS=4.3e-07 $X=79060 $Y=54745 $D=1
M196 546 49 306 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.4e-14 AS=1.15e-14 PD=4.8e-07 PS=4.3e-07 $X=79060 $Y=57825 $D=1
M197 GND CLK_MAIN 74 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.2e-14 AS=1.2e-14 PD=4.4e-07 PS=4.4e-07 $X=79410 $Y=49225 $D=1
M198 547 292 545 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.4e-14 AS=1.4e-14 PD=4.8e-07 PS=4.8e-07 $X=79440 $Y=54745 $D=1
M199 548 292 546 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.4e-14 AS=1.4e-14 PD=4.8e-07 PS=4.8e-07 $X=79440 $Y=57825 $D=1
M200 GND 84 295 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.2e-14 AS=1.2e-14 PD=4.4e-07 PS=4.4e-07 $X=79550 $Y=62980 $D=1
M201 GND 84 83 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.2e-14 AS=1.2e-14 PD=4.4e-07 PS=4.4e-07 $X=79550 $Y=63840 $D=1
M202 549 83 84 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.5e-14 AS=1.2e-14 PD=5e-07 PS=4.4e-07 $X=79550 $Y=64700 $D=1
M203 550 81 549 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.4e-14 AS=1.5e-14 PD=4.8e-07 PS=5e-07 $X=79550 $Y=65100 $D=1
M204 GND 80 550 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.2e-14 AS=1.4e-14 PD=4.4e-07 PS=4.8e-07 $X=79550 $Y=65480 $D=1
M205 GND RESET 81 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.2e-14 AS=1.2e-14 PD=4.4e-07 PS=4.4e-07 $X=79550 $Y=66360 $D=1
M206 GND 80 79 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.2e-14 AS=1.2e-14 PD=4.4e-07 PS=4.4e-07 $X=79550 $Y=67220 $D=1
M207 GND CLK_MAIN 80 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.2e-14 AS=1.2e-14 PD=4.4e-07 PS=4.4e-07 $X=79550 $Y=68080 $D=1
M208 85 79 84 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.2e-14 AS=1.2e-14 PD=4.4e-07 PS=4.4e-07 $X=79550 $Y=68940 $D=1
M209 551 79 GND GND NMOS_VTL L=5e-08 W=1e-07 AD=1.4e-14 AS=1.2e-14 PD=4.8e-07 PS=4.4e-07 $X=79550 $Y=69800 $D=1
M210 82 85 551 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.2e-14 AS=1.4e-14 PD=4.4e-07 PS=4.8e-07 $X=79550 $Y=70180 $D=1
M211 552 81 85 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.5e-14 AS=1.2e-14 PD=5e-07 PS=4.4e-07 $X=79550 $Y=71040 $D=1
M212 GND 82 552 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.2e-14 AS=1.5e-14 PD=4.4e-07 PS=5e-07 $X=79550 $Y=71440 $D=1
M213 307 80 82 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.2e-14 AS=1.2e-14 PD=4.4e-07 PS=4.4e-07 $X=79550 $Y=72300 $D=1
M214 GND 308 307 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.2e-14 AS=1.2e-14 PD=4.4e-07 PS=4.4e-07 $X=79550 $Y=73160 $D=1
M215 GND B2 308 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.2e-14 AS=1.2e-14 PD=4.4e-07 PS=4.4e-07 $X=79550 $Y=74020 $D=1
M216 GND 295 547 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.15e-14 AS=1.4e-14 PD=4.3e-07 PS=4.8e-07 $X=79820 $Y=54745 $D=1
M217 GND 295 548 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.15e-14 AS=1.4e-14 PD=4.3e-07 PS=4.8e-07 $X=79820 $Y=57825 $D=1
M218 86 75 67 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.2e-14 AS=1.2e-14 PD=4.4e-07 PS=4.4e-07 $X=80270 $Y=49225 $D=1
M219 91 305 GND GND NMOS_VTL L=5e-08 W=1e-07 AD=1.2e-14 AS=1.2e-14 PD=4.4e-07 PS=4.4e-07 $X=80925 $Y=55295 $D=1
M220 310 GND GND GND NMOS_VTL L=5e-08 W=1e-07 AD=1.35e-14 AS=1.15e-14 PD=4.7e-07 PS=4.3e-07 $X=80950 $Y=57465 $D=1
M221 553 75 GND GND NMOS_VTL L=5e-08 W=1e-07 AD=1.4e-14 AS=1.2e-14 PD=4.8e-07 PS=4.4e-07 $X=81130 $Y=49225 $D=1
M222 89 86 553 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.2e-14 AS=1.4e-14 PD=4.4e-07 PS=4.8e-07 $X=81510 $Y=49225 $D=1
M223 SC2 310 88 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.4e-14 AS=1.2e-14 PD=4.8e-07 PS=4.4e-07 $X=81720 $Y=57465 $D=1
M224 GND 306 88 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.2e-14 AS=1.2e-14 PD=4.4e-07 PS=4.4e-07 $X=81930 $Y=58615 $D=1
M225 91 GND SC2 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.15e-14 AS=1.4e-14 PD=4.3e-07 PS=4.8e-07 $X=82100 $Y=57465 $D=1
M226 554 76 86 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.5e-14 AS=1.2e-14 PD=5e-07 PS=4.4e-07 $X=82370 $Y=49225 $D=1
M227 GND 89 554 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.2e-14 AS=1.5e-14 PD=4.4e-07 PS=5e-07 $X=82770 $Y=49225 $D=1
M228 311 74 89 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.2e-14 AS=1.2e-14 PD=4.4e-07 PS=4.4e-07 $X=83630 $Y=49225 $D=1
M229 GND 312 311 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.2e-14 AS=1.2e-14 PD=4.4e-07 PS=4.4e-07 $X=84490 $Y=49225 $D=1
M230 GND SC2 312 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.2e-14 AS=1.2e-14 PD=4.4e-07 PS=4.4e-07 $X=85350 $Y=49225 $D=1
M231 GND 315 313 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.2e-14 AS=1.2e-14 PD=4.4e-07 PS=4.4e-07 $X=85755 $Y=61795 $D=1
M232 GND 97 315 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.2e-14 AS=1.2e-14 PD=4.4e-07 PS=4.4e-07 $X=85755 $Y=62980 $D=1
M233 GND 97 96 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.2e-14 AS=1.2e-14 PD=4.4e-07 PS=4.4e-07 $X=85755 $Y=63840 $D=1
M234 555 96 97 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.5e-14 AS=1.2e-14 PD=5e-07 PS=4.4e-07 $X=85755 $Y=64700 $D=1
M235 556 94 555 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.4e-14 AS=1.5e-14 PD=4.8e-07 PS=5e-07 $X=85755 $Y=65100 $D=1
M236 GND 93 556 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.2e-14 AS=1.4e-14 PD=4.4e-07 PS=4.8e-07 $X=85755 $Y=65480 $D=1
M237 GND RESET 94 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.2e-14 AS=1.2e-14 PD=4.4e-07 PS=4.4e-07 $X=85755 $Y=66360 $D=1
M238 GND 93 92 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.2e-14 AS=1.2e-14 PD=4.4e-07 PS=4.4e-07 $X=85755 $Y=67220 $D=1
M239 GND CLK_MAIN 93 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.2e-14 AS=1.2e-14 PD=4.4e-07 PS=4.4e-07 $X=85755 $Y=68080 $D=1
M240 98 92 97 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.2e-14 AS=1.2e-14 PD=4.4e-07 PS=4.4e-07 $X=85755 $Y=68940 $D=1
M241 557 92 GND GND NMOS_VTL L=5e-08 W=1e-07 AD=1.4e-14 AS=1.2e-14 PD=4.8e-07 PS=4.4e-07 $X=85755 $Y=69800 $D=1
M242 95 98 557 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.2e-14 AS=1.4e-14 PD=4.4e-07 PS=4.8e-07 $X=85755 $Y=70180 $D=1
M243 558 94 98 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.5e-14 AS=1.2e-14 PD=5e-07 PS=4.4e-07 $X=85755 $Y=71040 $D=1
M244 GND 95 558 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.2e-14 AS=1.5e-14 PD=4.4e-07 PS=5e-07 $X=85755 $Y=71440 $D=1
M245 316 93 95 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.2e-14 AS=1.2e-14 PD=4.4e-07 PS=4.4e-07 $X=85755 $Y=72300 $D=1
M246 GND 317 316 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.2e-14 AS=1.2e-14 PD=4.4e-07 PS=4.4e-07 $X=85755 $Y=73160 $D=1
M247 GND A3 317 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.2e-14 AS=1.2e-14 PD=4.4e-07 PS=4.4e-07 $X=85755 $Y=74020 $D=1
M248 GND 313 319 GND NMOS_VTL L=5e-08 W=1.15e-07 AD=1.61e-14 AS=1.3225e-14 PD=5.1e-07 PS=4.6e-07 $X=86390 $Y=54555 $D=1
M249 GND 313 321 GND NMOS_VTL L=5e-08 W=1.15e-07 AD=1.61e-14 AS=1.3225e-14 PD=5.1e-07 PS=4.6e-07 $X=86390 $Y=57635 $D=1
M250 GND 99 S3 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.2e-14 AS=1.2e-14 PD=4.4e-07 PS=4.4e-07 $X=86575 $Y=49225 $D=1
M251 319 318 GND GND NMOS_VTL L=5e-08 W=1.15e-07 AD=1.61e-14 AS=1.61e-14 PD=5.1e-07 PS=5.1e-07 $X=86770 $Y=54555 $D=1
M252 321 318 GND GND NMOS_VTL L=5e-08 W=1.15e-07 AD=1.61e-14 AS=1.61e-14 PD=5.1e-07 PS=5.1e-07 $X=86770 $Y=57635 $D=1
M253 106 77 319 GND NMOS_VTL L=5e-08 W=1.15e-07 AD=1.61e-14 AS=1.61e-14 PD=5.1e-07 PS=5.1e-07 $X=87150 $Y=54555 $D=1
M254 107 78 321 GND NMOS_VTL L=5e-08 W=1.15e-07 AD=1.61e-14 AS=1.61e-14 PD=5.1e-07 PS=5.1e-07 $X=87150 $Y=57635 $D=1
M255 GND 99 101 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.2e-14 AS=1.2e-14 PD=4.4e-07 PS=4.4e-07 $X=87435 $Y=49225 $D=1
M256 559 313 106 GND NMOS_VTL L=5e-08 W=1.15e-07 AD=1.61e-14 AS=1.61e-14 PD=5.1e-07 PS=5.1e-07 $X=87530 $Y=54555 $D=1
M257 560 313 107 GND NMOS_VTL L=5e-08 W=1.15e-07 AD=1.61e-14 AS=1.61e-14 PD=5.1e-07 PS=5.1e-07 $X=87530 $Y=57635 $D=1
M258 GND 318 559 GND NMOS_VTL L=5e-08 W=1.15e-07 AD=1.3225e-14 AS=1.61e-14 PD=4.6e-07 PS=5.1e-07 $X=87910 $Y=54555 $D=1
M259 GND 318 560 GND NMOS_VTL L=5e-08 W=1.15e-07 AD=1.3225e-14 AS=1.61e-14 PD=4.6e-07 PS=5.1e-07 $X=87910 $Y=57635 $D=1
M260 561 101 99 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.5e-14 AS=1.2e-14 PD=5e-07 PS=4.4e-07 $X=88295 $Y=49225 $D=1
M261 324 313 GND GND NMOS_VTL L=5e-08 W=1e-07 AD=1.4e-14 AS=1.15e-14 PD=4.8e-07 PS=4.3e-07 $X=88630 $Y=54585 $D=1
M262 326 313 GND GND NMOS_VTL L=5e-08 W=1e-07 AD=1.4e-14 AS=1.15e-14 PD=4.8e-07 PS=4.3e-07 $X=88630 $Y=57665 $D=1
M263 562 105 561 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.4e-14 AS=1.5e-14 PD=4.8e-07 PS=5e-07 $X=88695 $Y=49225 $D=1
M264 GND 318 324 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.4e-14 AS=1.4e-14 PD=4.8e-07 PS=4.8e-07 $X=89010 $Y=54585 $D=1
M265 GND 318 326 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.4e-14 AS=1.4e-14 PD=4.8e-07 PS=4.8e-07 $X=89010 $Y=57665 $D=1
M266 GND 103 562 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.2e-14 AS=1.4e-14 PD=4.4e-07 PS=4.8e-07 $X=89075 $Y=49225 $D=1
M267 324 77 GND GND NMOS_VTL L=5e-08 W=1e-07 AD=1.15e-14 AS=1.4e-14 PD=4.3e-07 PS=4.8e-07 $X=89390 $Y=54585 $D=1
M268 326 78 GND GND NMOS_VTL L=5e-08 W=1e-07 AD=1.15e-14 AS=1.4e-14 PD=4.3e-07 PS=4.8e-07 $X=89390 $Y=57665 $D=1
M269 GND RESET 105 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.2e-14 AS=1.2e-14 PD=4.4e-07 PS=4.4e-07 $X=89955 $Y=49225 $D=1
M270 120 106 324 GND NMOS_VTL L=5e-08 W=9e-08 AD=1.08e-14 AS=1.125e-14 PD=4.2e-07 PS=4.3e-07 $X=90130 $Y=54585 $D=1
M271 117 107 326 GND NMOS_VTL L=5e-08 W=9e-08 AD=1.08e-14 AS=1.125e-14 PD=4.2e-07 PS=4.3e-07 $X=90130 $Y=57665 $D=1
M272 GND 103 104 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.2e-14 AS=1.2e-14 PD=4.4e-07 PS=4.4e-07 $X=90815 $Y=49225 $D=1
M273 563 77 120 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.4e-14 AS=1.15e-14 PD=4.8e-07 PS=4.3e-07 $X=90860 $Y=54585 $D=1
M274 564 78 117 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.4e-14 AS=1.15e-14 PD=4.8e-07 PS=4.3e-07 $X=90860 $Y=57665 $D=1
M275 569 313 563 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.4e-14 AS=1.4e-14 PD=4.8e-07 PS=4.8e-07 $X=91240 $Y=54585 $D=1
M276 570 313 564 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.4e-14 AS=1.4e-14 PD=4.8e-07 PS=4.8e-07 $X=91240 $Y=57665 $D=1
M277 GND 328 318 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.2e-14 AS=1.2e-14 PD=4.4e-07 PS=4.4e-07 $X=91275 $Y=61795 $D=1
M278 GND 113 328 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.2e-14 AS=1.2e-14 PD=4.4e-07 PS=4.4e-07 $X=91275 $Y=62980 $D=1
M279 GND 113 112 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.2e-14 AS=1.2e-14 PD=4.4e-07 PS=4.4e-07 $X=91275 $Y=63840 $D=1
M280 565 112 113 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.5e-14 AS=1.2e-14 PD=5e-07 PS=4.4e-07 $X=91275 $Y=64700 $D=1
M281 566 110 565 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.4e-14 AS=1.5e-14 PD=4.8e-07 PS=5e-07 $X=91275 $Y=65100 $D=1
M282 GND 109 566 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.2e-14 AS=1.4e-14 PD=4.4e-07 PS=4.8e-07 $X=91275 $Y=65480 $D=1
M283 GND RESET 110 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.2e-14 AS=1.2e-14 PD=4.4e-07 PS=4.4e-07 $X=91275 $Y=66360 $D=1
M284 GND 109 108 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.2e-14 AS=1.2e-14 PD=4.4e-07 PS=4.4e-07 $X=91275 $Y=67220 $D=1
M285 GND CLK_MAIN 109 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.2e-14 AS=1.2e-14 PD=4.4e-07 PS=4.4e-07 $X=91275 $Y=68080 $D=1
M286 114 108 113 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.2e-14 AS=1.2e-14 PD=4.4e-07 PS=4.4e-07 $X=91275 $Y=68940 $D=1
M287 567 108 GND GND NMOS_VTL L=5e-08 W=1e-07 AD=1.4e-14 AS=1.2e-14 PD=4.8e-07 PS=4.4e-07 $X=91275 $Y=69800 $D=1
M288 111 114 567 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.2e-14 AS=1.4e-14 PD=4.4e-07 PS=4.8e-07 $X=91275 $Y=70180 $D=1
M289 568 110 114 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.5e-14 AS=1.2e-14 PD=5e-07 PS=4.4e-07 $X=91275 $Y=71040 $D=1
M290 GND 111 568 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.2e-14 AS=1.5e-14 PD=4.4e-07 PS=5e-07 $X=91275 $Y=71440 $D=1
M291 329 109 111 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.2e-14 AS=1.2e-14 PD=4.4e-07 PS=4.4e-07 $X=91275 $Y=72300 $D=1
M292 GND 330 329 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.2e-14 AS=1.2e-14 PD=4.4e-07 PS=4.4e-07 $X=91275 $Y=73160 $D=1
M293 GND B3 330 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.2e-14 AS=1.2e-14 PD=4.4e-07 PS=4.4e-07 $X=91275 $Y=74020 $D=1
M294 GND 318 569 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.15e-14 AS=1.4e-14 PD=4.3e-07 PS=4.8e-07 $X=91620 $Y=54585 $D=1
M295 GND 318 570 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.15e-14 AS=1.4e-14 PD=4.3e-07 PS=4.8e-07 $X=91620 $Y=57665 $D=1
M296 GND CLK_MAIN 103 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.2e-14 AS=1.2e-14 PD=4.4e-07 PS=4.4e-07 $X=91675 $Y=49225 $D=1
M297 116 104 99 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.2e-14 AS=1.2e-14 PD=4.4e-07 PS=4.4e-07 $X=92535 $Y=49225 $D=1
M298 332 GND GND GND NMOS_VTL L=5e-08 W=1e-07 AD=1.35e-14 AS=1.15e-14 PD=4.7e-07 PS=4.3e-07 $X=92750 $Y=57305 $D=1
M299 571 104 GND GND NMOS_VTL L=5e-08 W=1e-07 AD=1.4e-14 AS=1.2e-14 PD=4.8e-07 PS=4.4e-07 $X=93395 $Y=49225 $D=1
M300 SC3 332 117 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.4e-14 AS=1.2e-14 PD=4.8e-07 PS=4.4e-07 $X=93520 $Y=57305 $D=1
M301 119 116 571 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.2e-14 AS=1.4e-14 PD=4.4e-07 PS=4.8e-07 $X=93775 $Y=49225 $D=1
M302 120 GND SC3 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.15e-14 AS=1.4e-14 PD=4.3e-07 PS=4.8e-07 $X=93900 $Y=57305 $D=1
M303 572 105 116 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.5e-14 AS=1.2e-14 PD=5e-07 PS=4.4e-07 $X=94635 $Y=49225 $D=1
M304 GND 119 572 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.2e-14 AS=1.5e-14 PD=4.4e-07 PS=5e-07 $X=95035 $Y=49225 $D=1
M305 333 GND GND GND NMOS_VTL L=5e-08 W=1e-07 AD=1.35e-14 AS=1.15e-14 PD=4.7e-07 PS=4.3e-07 $X=95855 $Y=57280 $D=1
M306 334 103 119 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.2e-14 AS=1.2e-14 PD=4.4e-07 PS=4.4e-07 $X=95895 $Y=49225 $D=1
M307 121 333 107 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.4e-14 AS=1.2e-14 PD=4.8e-07 PS=4.4e-07 $X=96625 $Y=57280 $D=1
M308 GND 335 334 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.2e-14 AS=1.2e-14 PD=4.4e-07 PS=4.4e-07 $X=96755 $Y=49225 $D=1
M309 106 GND 121 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.15e-14 AS=1.4e-14 PD=4.3e-07 PS=4.8e-07 $X=97005 $Y=57280 $D=1
M310 GND SC3 335 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.2e-14 AS=1.2e-14 PD=4.4e-07 PS=4.4e-07 $X=97615 $Y=49225 $D=1
M311 GND 122 S4 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.2e-14 AS=1.2e-14 PD=4.4e-07 PS=4.4e-07 $X=99550 $Y=49225 $D=1
M312 GND 122 123 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.2e-14 AS=1.2e-14 PD=4.4e-07 PS=4.4e-07 $X=100410 $Y=49225 $D=1
M313 GND 130 337 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.2e-14 AS=1.2e-14 PD=4.4e-07 PS=4.4e-07 $X=100920 $Y=62980 $D=1
M314 GND 130 129 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.2e-14 AS=1.2e-14 PD=4.4e-07 PS=4.4e-07 $X=100920 $Y=63840 $D=1
M315 573 129 130 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.5e-14 AS=1.2e-14 PD=5e-07 PS=4.4e-07 $X=100920 $Y=64700 $D=1
M316 574 127 573 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.4e-14 AS=1.5e-14 PD=4.8e-07 PS=5e-07 $X=100920 $Y=65100 $D=1
M317 GND 125 574 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.2e-14 AS=1.4e-14 PD=4.4e-07 PS=4.8e-07 $X=100920 $Y=65480 $D=1
M318 GND RESET 127 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.2e-14 AS=1.2e-14 PD=4.4e-07 PS=4.4e-07 $X=100920 $Y=66360 $D=1
M319 GND 125 124 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.2e-14 AS=1.2e-14 PD=4.4e-07 PS=4.4e-07 $X=100920 $Y=67220 $D=1
M320 GND CLK_MAIN 125 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.2e-14 AS=1.2e-14 PD=4.4e-07 PS=4.4e-07 $X=100920 $Y=68080 $D=1
M321 131 124 130 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.2e-14 AS=1.2e-14 PD=4.4e-07 PS=4.4e-07 $X=100920 $Y=68940 $D=1
M322 575 124 GND GND NMOS_VTL L=5e-08 W=1e-07 AD=1.4e-14 AS=1.2e-14 PD=4.8e-07 PS=4.4e-07 $X=100920 $Y=69800 $D=1
M323 128 131 575 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.2e-14 AS=1.4e-14 PD=4.4e-07 PS=4.8e-07 $X=100920 $Y=70180 $D=1
M324 576 127 131 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.5e-14 AS=1.2e-14 PD=5e-07 PS=4.4e-07 $X=100920 $Y=71040 $D=1
M325 GND 128 576 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.2e-14 AS=1.5e-14 PD=4.4e-07 PS=5e-07 $X=100920 $Y=71440 $D=1
M326 338 125 128 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.2e-14 AS=1.2e-14 PD=4.4e-07 PS=4.4e-07 $X=100920 $Y=72300 $D=1
M327 GND 339 338 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.2e-14 AS=1.2e-14 PD=4.4e-07 PS=4.4e-07 $X=100920 $Y=73160 $D=1
M328 GND A4 339 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.2e-14 AS=1.2e-14 PD=4.4e-07 PS=4.4e-07 $X=100920 $Y=74020 $D=1
M329 577 123 122 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.5e-14 AS=1.2e-14 PD=5e-07 PS=4.4e-07 $X=101270 $Y=49225 $D=1
M330 GND 337 341 GND NMOS_VTL L=5e-08 W=1.15e-07 AD=1.61e-14 AS=1.3225e-14 PD=5.1e-07 PS=4.6e-07 $X=101460 $Y=54715 $D=1
M331 GND 337 343 GND NMOS_VTL L=5e-08 W=1.15e-07 AD=1.61e-14 AS=1.3225e-14 PD=5.1e-07 PS=4.6e-07 $X=101460 $Y=57635 $D=1
M332 578 135 577 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.4e-14 AS=1.5e-14 PD=4.8e-07 PS=5e-07 $X=101670 $Y=49225 $D=1
M333 341 340 GND GND NMOS_VTL L=5e-08 W=1.15e-07 AD=1.61e-14 AS=1.61e-14 PD=5.1e-07 PS=5.1e-07 $X=101840 $Y=54715 $D=1
M334 343 340 GND GND NMOS_VTL L=5e-08 W=1.15e-07 AD=1.61e-14 AS=1.61e-14 PD=5.1e-07 PS=5.1e-07 $X=101840 $Y=57635 $D=1
M335 GND 133 578 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.2e-14 AS=1.4e-14 PD=4.4e-07 PS=4.8e-07 $X=102050 $Y=49225 $D=1
M336 136 VDD 341 GND NMOS_VTL L=5e-08 W=1.15e-07 AD=1.61e-14 AS=1.61e-14 PD=5.1e-07 PS=5.1e-07 $X=102220 $Y=54715 $D=1
M337 137 GND 343 GND NMOS_VTL L=5e-08 W=1.15e-07 AD=1.61e-14 AS=1.61e-14 PD=5.1e-07 PS=5.1e-07 $X=102220 $Y=57635 $D=1
M338 579 337 136 GND NMOS_VTL L=5e-08 W=1.15e-07 AD=1.61e-14 AS=1.61e-14 PD=5.1e-07 PS=5.1e-07 $X=102600 $Y=54715 $D=1
M339 580 337 137 GND NMOS_VTL L=5e-08 W=1.15e-07 AD=1.61e-14 AS=1.61e-14 PD=5.1e-07 PS=5.1e-07 $X=102600 $Y=57635 $D=1
M340 GND RESET 135 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.2e-14 AS=1.2e-14 PD=4.4e-07 PS=4.4e-07 $X=102930 $Y=49225 $D=1
M341 GND 340 579 GND NMOS_VTL L=5e-08 W=1.15e-07 AD=1.3225e-14 AS=1.61e-14 PD=4.6e-07 PS=5.1e-07 $X=102980 $Y=54715 $D=1
M342 GND 340 580 GND NMOS_VTL L=5e-08 W=1.15e-07 AD=1.3225e-14 AS=1.61e-14 PD=4.6e-07 PS=5.1e-07 $X=102980 $Y=57635 $D=1
M343 346 337 GND GND NMOS_VTL L=5e-08 W=1e-07 AD=1.4e-14 AS=1.15e-14 PD=4.8e-07 PS=4.3e-07 $X=103700 $Y=54745 $D=1
M344 348 337 GND GND NMOS_VTL L=5e-08 W=1e-07 AD=1.4e-14 AS=1.15e-14 PD=4.8e-07 PS=4.3e-07 $X=103700 $Y=57665 $D=1
M345 GND 133 134 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.2e-14 AS=1.2e-14 PD=4.4e-07 PS=4.4e-07 $X=103790 $Y=49225 $D=1
M346 GND 340 346 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.4e-14 AS=1.4e-14 PD=4.8e-07 PS=4.8e-07 $X=104080 $Y=54745 $D=1
M347 GND 340 348 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.4e-14 AS=1.4e-14 PD=4.8e-07 PS=4.8e-07 $X=104080 $Y=57665 $D=1
M348 346 VDD GND GND NMOS_VTL L=5e-08 W=1e-07 AD=1.15e-14 AS=1.4e-14 PD=4.3e-07 PS=4.8e-07 $X=104460 $Y=54745 $D=1
M349 348 GND GND GND NMOS_VTL L=5e-08 W=1e-07 AD=1.15e-14 AS=1.4e-14 PD=4.3e-07 PS=4.8e-07 $X=104460 $Y=57665 $D=1
M350 GND CLK_MAIN 133 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.2e-14 AS=1.2e-14 PD=4.4e-07 PS=4.4e-07 $X=104650 $Y=49225 $D=1
M351 350 136 346 GND NMOS_VTL L=5e-08 W=9e-08 AD=1.08e-14 AS=1.125e-14 PD=4.2e-07 PS=4.3e-07 $X=105200 $Y=54745 $D=1
M352 351 137 348 GND NMOS_VTL L=5e-08 W=9e-08 AD=1.08e-14 AS=1.125e-14 PD=4.2e-07 PS=4.3e-07 $X=105200 $Y=57665 $D=1
M353 139 134 122 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.2e-14 AS=1.2e-14 PD=4.4e-07 PS=4.4e-07 $X=105510 $Y=49225 $D=1
M354 581 VDD 350 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.4e-14 AS=1.15e-14 PD=4.8e-07 PS=4.3e-07 $X=105930 $Y=54745 $D=1
M355 582 GND 351 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.4e-14 AS=1.15e-14 PD=4.8e-07 PS=4.3e-07 $X=105930 $Y=57665 $D=1
M356 583 337 581 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.4e-14 AS=1.4e-14 PD=4.8e-07 PS=4.8e-07 $X=106310 $Y=54745 $D=1
M357 584 337 582 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.4e-14 AS=1.4e-14 PD=4.8e-07 PS=4.8e-07 $X=106310 $Y=57665 $D=1
M358 589 134 GND GND NMOS_VTL L=5e-08 W=1e-07 AD=1.4e-14 AS=1.2e-14 PD=4.8e-07 PS=4.4e-07 $X=106370 $Y=49225 $D=1
M359 GND 144 340 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.2e-14 AS=1.2e-14 PD=4.4e-07 PS=4.4e-07 $X=106420 $Y=62980 $D=1
M360 GND 144 143 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.2e-14 AS=1.2e-14 PD=4.4e-07 PS=4.4e-07 $X=106420 $Y=63840 $D=1
M361 585 143 144 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.5e-14 AS=1.2e-14 PD=5e-07 PS=4.4e-07 $X=106420 $Y=64700 $D=1
M362 586 141 585 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.4e-14 AS=1.5e-14 PD=4.8e-07 PS=5e-07 $X=106420 $Y=65100 $D=1
M363 GND 140 586 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.2e-14 AS=1.4e-14 PD=4.4e-07 PS=4.8e-07 $X=106420 $Y=65480 $D=1
M364 GND RESET 141 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.2e-14 AS=1.2e-14 PD=4.4e-07 PS=4.4e-07 $X=106420 $Y=66360 $D=1
M365 GND 140 138 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.2e-14 AS=1.2e-14 PD=4.4e-07 PS=4.4e-07 $X=106420 $Y=67220 $D=1
M366 GND CLK_MAIN 140 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.2e-14 AS=1.2e-14 PD=4.4e-07 PS=4.4e-07 $X=106420 $Y=68080 $D=1
M367 145 138 144 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.2e-14 AS=1.2e-14 PD=4.4e-07 PS=4.4e-07 $X=106420 $Y=68940 $D=1
M368 587 138 GND GND NMOS_VTL L=5e-08 W=1e-07 AD=1.4e-14 AS=1.2e-14 PD=4.8e-07 PS=4.4e-07 $X=106420 $Y=69800 $D=1
M369 142 145 587 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.2e-14 AS=1.4e-14 PD=4.4e-07 PS=4.8e-07 $X=106420 $Y=70180 $D=1
M370 588 141 145 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.5e-14 AS=1.2e-14 PD=5e-07 PS=4.4e-07 $X=106420 $Y=71040 $D=1
M371 GND 142 588 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.2e-14 AS=1.5e-14 PD=4.4e-07 PS=5e-07 $X=106420 $Y=71440 $D=1
M372 352 140 142 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.2e-14 AS=1.2e-14 PD=4.4e-07 PS=4.4e-07 $X=106420 $Y=72300 $D=1
M373 GND 353 352 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.2e-14 AS=1.2e-14 PD=4.4e-07 PS=4.4e-07 $X=106420 $Y=73160 $D=1
M374 GND B4 353 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.2e-14 AS=1.2e-14 PD=4.4e-07 PS=4.4e-07 $X=106420 $Y=74020 $D=1
M375 GND 340 583 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.15e-14 AS=1.4e-14 PD=4.3e-07 PS=4.8e-07 $X=106690 $Y=54745 $D=1
M376 GND 340 584 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.15e-14 AS=1.4e-14 PD=4.3e-07 PS=4.8e-07 $X=106690 $Y=57665 $D=1
M377 146 139 589 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.2e-14 AS=1.4e-14 PD=4.4e-07 PS=4.8e-07 $X=106750 $Y=49225 $D=1
M378 590 135 139 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.5e-14 AS=1.2e-14 PD=5e-07 PS=4.4e-07 $X=107610 $Y=49225 $D=1
M379 150 350 GND GND NMOS_VTL L=5e-08 W=1e-07 AD=1.2e-14 AS=1.2e-14 PD=4.4e-07 PS=4.4e-07 $X=107795 $Y=55295 $D=1
M380 355 121 GND GND NMOS_VTL L=5e-08 W=1e-07 AD=1.35e-14 AS=1.15e-14 PD=4.7e-07 PS=4.3e-07 $X=107820 $Y=57305 $D=1
M381 GND 146 590 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.2e-14 AS=1.5e-14 PD=4.4e-07 PS=5e-07 $X=108010 $Y=49225 $D=1
M382 SC4 355 148 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.4e-14 AS=1.2e-14 PD=4.8e-07 PS=4.4e-07 $X=108590 $Y=57305 $D=1
M383 GND 351 148 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.2e-14 AS=1.2e-14 PD=4.4e-07 PS=4.4e-07 $X=108800 $Y=58455 $D=1
M384 356 133 146 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.2e-14 AS=1.2e-14 PD=4.4e-07 PS=4.4e-07 $X=108870 $Y=49225 $D=1
M385 150 121 SC4 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.15e-14 AS=1.4e-14 PD=4.3e-07 PS=4.8e-07 $X=108970 $Y=57305 $D=1
M386 GND 357 356 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.2e-14 AS=1.2e-14 PD=4.4e-07 PS=4.4e-07 $X=109730 $Y=49225 $D=1
M387 GND SC4 357 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.2e-14 AS=1.2e-14 PD=4.4e-07 PS=4.4e-07 $X=110590 $Y=49225 $D=1
M388 GND 153 S5 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.2e-14 AS=1.2e-14 PD=4.4e-07 PS=4.4e-07 $X=111970 $Y=49225 $D=1
M389 GND 360 359 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.2e-14 AS=1.2e-14 PD=4.4e-07 PS=4.4e-07 $X=112625 $Y=61795 $D=1
M390 GND 158 360 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.2e-14 AS=1.2e-14 PD=4.4e-07 PS=4.4e-07 $X=112625 $Y=62980 $D=1
M391 GND 158 157 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.2e-14 AS=1.2e-14 PD=4.4e-07 PS=4.4e-07 $X=112625 $Y=63840 $D=1
M392 591 157 158 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.5e-14 AS=1.2e-14 PD=5e-07 PS=4.4e-07 $X=112625 $Y=64700 $D=1
M393 592 155 591 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.4e-14 AS=1.5e-14 PD=4.8e-07 PS=5e-07 $X=112625 $Y=65100 $D=1
M394 GND 152 592 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.2e-14 AS=1.4e-14 PD=4.4e-07 PS=4.8e-07 $X=112625 $Y=65480 $D=1
M395 GND RESET 155 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.2e-14 AS=1.2e-14 PD=4.4e-07 PS=4.4e-07 $X=112625 $Y=66360 $D=1
M396 GND 152 151 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.2e-14 AS=1.2e-14 PD=4.4e-07 PS=4.4e-07 $X=112625 $Y=67220 $D=1
M397 GND CLK_MAIN 152 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.2e-14 AS=1.2e-14 PD=4.4e-07 PS=4.4e-07 $X=112625 $Y=68080 $D=1
M398 159 151 158 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.2e-14 AS=1.2e-14 PD=4.4e-07 PS=4.4e-07 $X=112625 $Y=68940 $D=1
M399 593 151 GND GND NMOS_VTL L=5e-08 W=1e-07 AD=1.4e-14 AS=1.2e-14 PD=4.8e-07 PS=4.4e-07 $X=112625 $Y=69800 $D=1
M400 156 159 593 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.2e-14 AS=1.4e-14 PD=4.4e-07 PS=4.8e-07 $X=112625 $Y=70180 $D=1
M401 594 155 159 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.5e-14 AS=1.2e-14 PD=5e-07 PS=4.4e-07 $X=112625 $Y=71040 $D=1
M402 GND 156 594 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.2e-14 AS=1.5e-14 PD=4.4e-07 PS=5e-07 $X=112625 $Y=71440 $D=1
M403 361 152 156 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.2e-14 AS=1.2e-14 PD=4.4e-07 PS=4.4e-07 $X=112625 $Y=72300 $D=1
M404 GND 362 361 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.2e-14 AS=1.2e-14 PD=4.4e-07 PS=4.4e-07 $X=112625 $Y=73160 $D=1
M405 GND A5 362 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.2e-14 AS=1.2e-14 PD=4.4e-07 PS=4.4e-07 $X=112625 $Y=74020 $D=1
M406 GND 153 154 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.2e-14 AS=1.2e-14 PD=4.4e-07 PS=4.4e-07 $X=112830 $Y=49225 $D=1
M407 GND 359 364 GND NMOS_VTL L=5e-08 W=1.15e-07 AD=1.61e-14 AS=1.3225e-14 PD=5.1e-07 PS=4.6e-07 $X=113260 $Y=54505 $D=1
M408 GND 359 366 GND NMOS_VTL L=5e-08 W=1.15e-07 AD=1.61e-14 AS=1.3225e-14 PD=5.1e-07 PS=4.6e-07 $X=113260 $Y=57585 $D=1
M409 364 363 GND GND NMOS_VTL L=5e-08 W=1.15e-07 AD=1.61e-14 AS=1.61e-14 PD=5.1e-07 PS=5.1e-07 $X=113640 $Y=54505 $D=1
M410 366 363 GND GND NMOS_VTL L=5e-08 W=1.15e-07 AD=1.61e-14 AS=1.61e-14 PD=5.1e-07 PS=5.1e-07 $X=113640 $Y=57585 $D=1
M411 595 154 153 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.5e-14 AS=1.2e-14 PD=5e-07 PS=4.4e-07 $X=113690 $Y=49225 $D=1
M412 165 136 364 GND NMOS_VTL L=5e-08 W=1.15e-07 AD=1.61e-14 AS=1.61e-14 PD=5.1e-07 PS=5.1e-07 $X=114020 $Y=54505 $D=1
M413 166 137 366 GND NMOS_VTL L=5e-08 W=1.15e-07 AD=1.61e-14 AS=1.61e-14 PD=5.1e-07 PS=5.1e-07 $X=114020 $Y=57585 $D=1
M414 596 164 595 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.4e-14 AS=1.5e-14 PD=4.8e-07 PS=5e-07 $X=114090 $Y=49225 $D=1
M415 597 359 165 GND NMOS_VTL L=5e-08 W=1.15e-07 AD=1.61e-14 AS=1.61e-14 PD=5.1e-07 PS=5.1e-07 $X=114400 $Y=54505 $D=1
M416 598 359 166 GND NMOS_VTL L=5e-08 W=1.15e-07 AD=1.61e-14 AS=1.61e-14 PD=5.1e-07 PS=5.1e-07 $X=114400 $Y=57585 $D=1
M417 GND 162 596 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.2e-14 AS=1.4e-14 PD=4.4e-07 PS=4.8e-07 $X=114470 $Y=49225 $D=1
M418 GND 363 597 GND NMOS_VTL L=5e-08 W=1.15e-07 AD=1.3225e-14 AS=1.61e-14 PD=4.6e-07 PS=5.1e-07 $X=114780 $Y=54505 $D=1
M419 GND 363 598 GND NMOS_VTL L=5e-08 W=1.15e-07 AD=1.3225e-14 AS=1.61e-14 PD=4.6e-07 PS=5.1e-07 $X=114780 $Y=57585 $D=1
M420 GND RESET 164 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.2e-14 AS=1.2e-14 PD=4.4e-07 PS=4.4e-07 $X=115350 $Y=49225 $D=1
M421 369 359 GND GND NMOS_VTL L=5e-08 W=1e-07 AD=1.4e-14 AS=1.15e-14 PD=4.8e-07 PS=4.3e-07 $X=115500 $Y=54535 $D=1
M422 371 359 GND GND NMOS_VTL L=5e-08 W=1e-07 AD=1.4e-14 AS=1.15e-14 PD=4.8e-07 PS=4.3e-07 $X=115500 $Y=57615 $D=1
M423 GND 363 369 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.4e-14 AS=1.4e-14 PD=4.8e-07 PS=4.8e-07 $X=115880 $Y=54535 $D=1
M424 GND 363 371 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.4e-14 AS=1.4e-14 PD=4.8e-07 PS=4.8e-07 $X=115880 $Y=57615 $D=1
M425 GND 162 163 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.2e-14 AS=1.2e-14 PD=4.4e-07 PS=4.4e-07 $X=116210 $Y=49225 $D=1
M426 369 136 GND GND NMOS_VTL L=5e-08 W=1e-07 AD=1.15e-14 AS=1.4e-14 PD=4.3e-07 PS=4.8e-07 $X=116260 $Y=54535 $D=1
M427 371 137 GND GND NMOS_VTL L=5e-08 W=1e-07 AD=1.15e-14 AS=1.4e-14 PD=4.3e-07 PS=4.8e-07 $X=116260 $Y=57615 $D=1
M428 179 165 369 GND NMOS_VTL L=5e-08 W=9e-08 AD=1.08e-14 AS=1.125e-14 PD=4.2e-07 PS=4.3e-07 $X=117000 $Y=54535 $D=1
M429 177 166 371 GND NMOS_VTL L=5e-08 W=9e-08 AD=1.08e-14 AS=1.125e-14 PD=4.2e-07 PS=4.3e-07 $X=117000 $Y=57615 $D=1
M430 GND CLK_MAIN 162 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.2e-14 AS=1.2e-14 PD=4.4e-07 PS=4.4e-07 $X=117070 $Y=49225 $D=1
M431 599 136 179 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.4e-14 AS=1.15e-14 PD=4.8e-07 PS=4.3e-07 $X=117730 $Y=54535 $D=1
M432 600 137 177 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.4e-14 AS=1.15e-14 PD=4.8e-07 PS=4.3e-07 $X=117730 $Y=57615 $D=1
M433 169 163 153 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.2e-14 AS=1.2e-14 PD=4.4e-07 PS=4.4e-07 $X=117930 $Y=49225 $D=1
M434 605 359 599 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.4e-14 AS=1.4e-14 PD=4.8e-07 PS=4.8e-07 $X=118110 $Y=54535 $D=1
M435 606 359 600 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.4e-14 AS=1.4e-14 PD=4.8e-07 PS=4.8e-07 $X=118110 $Y=57615 $D=1
M436 GND 373 363 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.2e-14 AS=1.2e-14 PD=4.4e-07 PS=4.4e-07 $X=118145 $Y=61795 $D=1
M437 GND 173 373 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.2e-14 AS=1.2e-14 PD=4.4e-07 PS=4.4e-07 $X=118145 $Y=62980 $D=1
M438 GND 173 172 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.2e-14 AS=1.2e-14 PD=4.4e-07 PS=4.4e-07 $X=118145 $Y=63840 $D=1
M439 601 172 173 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.5e-14 AS=1.2e-14 PD=5e-07 PS=4.4e-07 $X=118145 $Y=64700 $D=1
M440 602 170 601 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.4e-14 AS=1.5e-14 PD=4.8e-07 PS=5e-07 $X=118145 $Y=65100 $D=1
M441 GND 168 602 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.2e-14 AS=1.4e-14 PD=4.4e-07 PS=4.8e-07 $X=118145 $Y=65480 $D=1
M442 GND RESET 170 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.2e-14 AS=1.2e-14 PD=4.4e-07 PS=4.4e-07 $X=118145 $Y=66360 $D=1
M443 GND 168 167 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.2e-14 AS=1.2e-14 PD=4.4e-07 PS=4.4e-07 $X=118145 $Y=67220 $D=1
M444 GND CLK_MAIN 168 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.2e-14 AS=1.2e-14 PD=4.4e-07 PS=4.4e-07 $X=118145 $Y=68080 $D=1
M445 174 167 173 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.2e-14 AS=1.2e-14 PD=4.4e-07 PS=4.4e-07 $X=118145 $Y=68940 $D=1
M446 603 167 GND GND NMOS_VTL L=5e-08 W=1e-07 AD=1.4e-14 AS=1.2e-14 PD=4.8e-07 PS=4.4e-07 $X=118145 $Y=69800 $D=1
M447 171 174 603 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.2e-14 AS=1.4e-14 PD=4.4e-07 PS=4.8e-07 $X=118145 $Y=70180 $D=1
M448 604 170 174 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.5e-14 AS=1.2e-14 PD=5e-07 PS=4.4e-07 $X=118145 $Y=71040 $D=1
M449 GND 171 604 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.2e-14 AS=1.5e-14 PD=4.4e-07 PS=5e-07 $X=118145 $Y=71440 $D=1
M450 374 168 171 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.2e-14 AS=1.2e-14 PD=4.4e-07 PS=4.4e-07 $X=118145 $Y=72300 $D=1
M451 GND 375 374 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.2e-14 AS=1.2e-14 PD=4.4e-07 PS=4.4e-07 $X=118145 $Y=73160 $D=1
M452 GND B5 375 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.2e-14 AS=1.2e-14 PD=4.4e-07 PS=4.4e-07 $X=118145 $Y=74020 $D=1
M453 GND 363 605 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.15e-14 AS=1.4e-14 PD=4.3e-07 PS=4.8e-07 $X=118490 $Y=54535 $D=1
M454 GND 363 606 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.15e-14 AS=1.4e-14 PD=4.3e-07 PS=4.8e-07 $X=118490 $Y=57615 $D=1
M455 607 163 GND GND NMOS_VTL L=5e-08 W=1e-07 AD=1.4e-14 AS=1.2e-14 PD=4.8e-07 PS=4.4e-07 $X=118790 $Y=49225 $D=1
M456 176 169 607 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.2e-14 AS=1.4e-14 PD=4.4e-07 PS=4.8e-07 $X=119170 $Y=49225 $D=1
M457 377 121 GND GND NMOS_VTL L=5e-08 W=1e-07 AD=1.35e-14 AS=1.15e-14 PD=4.7e-07 PS=4.3e-07 $X=119620 $Y=57255 $D=1
M458 608 164 169 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.5e-14 AS=1.2e-14 PD=5e-07 PS=4.4e-07 $X=120030 $Y=49225 $D=1
M459 SC5 377 177 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.4e-14 AS=1.2e-14 PD=4.8e-07 PS=4.4e-07 $X=120390 $Y=57255 $D=1
M460 GND 176 608 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.2e-14 AS=1.5e-14 PD=4.4e-07 PS=5e-07 $X=120430 $Y=49225 $D=1
M461 179 121 SC5 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.15e-14 AS=1.4e-14 PD=4.3e-07 PS=4.8e-07 $X=120770 $Y=57255 $D=1
M462 378 162 176 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.2e-14 AS=1.2e-14 PD=4.4e-07 PS=4.4e-07 $X=121290 $Y=49225 $D=1
M463 GND 379 378 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.2e-14 AS=1.2e-14 PD=4.4e-07 PS=4.4e-07 $X=122150 $Y=49225 $D=1
M464 GND SC5 379 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.2e-14 AS=1.2e-14 PD=4.4e-07 PS=4.4e-07 $X=123010 $Y=49225 $D=1
M465 GND 187 381 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.2e-14 AS=1.2e-14 PD=4.4e-07 PS=4.4e-07 $X=124520 $Y=62980 $D=1
M466 GND 187 186 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.2e-14 AS=1.2e-14 PD=4.4e-07 PS=4.4e-07 $X=124520 $Y=63840 $D=1
M467 609 186 187 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.5e-14 AS=1.2e-14 PD=5e-07 PS=4.4e-07 $X=124520 $Y=64700 $D=1
M468 610 183 609 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.4e-14 AS=1.5e-14 PD=4.8e-07 PS=5e-07 $X=124520 $Y=65100 $D=1
M469 GND 181 610 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.2e-14 AS=1.4e-14 PD=4.4e-07 PS=4.8e-07 $X=124520 $Y=65480 $D=1
M470 GND RESET 183 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.2e-14 AS=1.2e-14 PD=4.4e-07 PS=4.4e-07 $X=124520 $Y=66360 $D=1
M471 GND 181 180 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.2e-14 AS=1.2e-14 PD=4.4e-07 PS=4.4e-07 $X=124520 $Y=67220 $D=1
M472 GND CLK_MAIN 181 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.2e-14 AS=1.2e-14 PD=4.4e-07 PS=4.4e-07 $X=124520 $Y=68080 $D=1
M473 188 180 187 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.2e-14 AS=1.2e-14 PD=4.4e-07 PS=4.4e-07 $X=124520 $Y=68940 $D=1
M474 611 180 GND GND NMOS_VTL L=5e-08 W=1e-07 AD=1.4e-14 AS=1.2e-14 PD=4.8e-07 PS=4.4e-07 $X=124520 $Y=69800 $D=1
M475 184 188 611 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.2e-14 AS=1.4e-14 PD=4.4e-07 PS=4.8e-07 $X=124520 $Y=70180 $D=1
M476 612 183 188 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.5e-14 AS=1.2e-14 PD=5e-07 PS=4.4e-07 $X=124520 $Y=71040 $D=1
M477 GND 184 612 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.2e-14 AS=1.5e-14 PD=4.4e-07 PS=5e-07 $X=124520 $Y=71440 $D=1
M478 382 181 184 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.2e-14 AS=1.2e-14 PD=4.4e-07 PS=4.4e-07 $X=124520 $Y=72300 $D=1
M479 GND 383 382 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.2e-14 AS=1.2e-14 PD=4.4e-07 PS=4.4e-07 $X=124520 $Y=73160 $D=1
M480 GND A6 383 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.2e-14 AS=1.2e-14 PD=4.4e-07 PS=4.4e-07 $X=124520 $Y=74020 $D=1
M481 GND 182 S6 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.2e-14 AS=1.2e-14 PD=4.4e-07 PS=4.4e-07 $X=124525 $Y=49225 $D=1
M482 GND 381 385 GND NMOS_VTL L=5e-08 W=1.15e-07 AD=1.61e-14 AS=1.3225e-14 PD=5.1e-07 PS=4.6e-07 $X=125060 $Y=54555 $D=1
M483 GND 381 387 GND NMOS_VTL L=5e-08 W=1.15e-07 AD=1.61e-14 AS=1.3225e-14 PD=5.1e-07 PS=4.6e-07 $X=125060 $Y=57635 $D=1
M484 GND 182 185 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.2e-14 AS=1.2e-14 PD=4.4e-07 PS=4.4e-07 $X=125385 $Y=49225 $D=1
M485 385 384 GND GND NMOS_VTL L=5e-08 W=1.15e-07 AD=1.61e-14 AS=1.61e-14 PD=5.1e-07 PS=5.1e-07 $X=125440 $Y=54555 $D=1
M486 387 384 GND GND NMOS_VTL L=5e-08 W=1.15e-07 AD=1.61e-14 AS=1.61e-14 PD=5.1e-07 PS=5.1e-07 $X=125440 $Y=57635 $D=1
M487 194 165 385 GND NMOS_VTL L=5e-08 W=1.15e-07 AD=1.61e-14 AS=1.61e-14 PD=5.1e-07 PS=5.1e-07 $X=125820 $Y=54555 $D=1
M488 195 166 387 GND NMOS_VTL L=5e-08 W=1.15e-07 AD=1.61e-14 AS=1.61e-14 PD=5.1e-07 PS=5.1e-07 $X=125820 $Y=57635 $D=1
M489 613 381 194 GND NMOS_VTL L=5e-08 W=1.15e-07 AD=1.61e-14 AS=1.61e-14 PD=5.1e-07 PS=5.1e-07 $X=126200 $Y=54555 $D=1
M490 614 381 195 GND NMOS_VTL L=5e-08 W=1.15e-07 AD=1.61e-14 AS=1.61e-14 PD=5.1e-07 PS=5.1e-07 $X=126200 $Y=57635 $D=1
M491 615 185 182 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.5e-14 AS=1.2e-14 PD=5e-07 PS=4.4e-07 $X=126245 $Y=49225 $D=1
M492 GND 384 613 GND NMOS_VTL L=5e-08 W=1.15e-07 AD=1.3225e-14 AS=1.61e-14 PD=4.6e-07 PS=5.1e-07 $X=126580 $Y=54555 $D=1
M493 GND 384 614 GND NMOS_VTL L=5e-08 W=1.15e-07 AD=1.3225e-14 AS=1.61e-14 PD=4.6e-07 PS=5.1e-07 $X=126580 $Y=57635 $D=1
M494 616 193 615 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.4e-14 AS=1.5e-14 PD=4.8e-07 PS=5e-07 $X=126645 $Y=49225 $D=1
M495 GND 191 616 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.2e-14 AS=1.4e-14 PD=4.4e-07 PS=4.8e-07 $X=127025 $Y=49225 $D=1
M496 390 381 GND GND NMOS_VTL L=5e-08 W=1e-07 AD=1.4e-14 AS=1.15e-14 PD=4.8e-07 PS=4.3e-07 $X=127300 $Y=54585 $D=1
M497 392 381 GND GND NMOS_VTL L=5e-08 W=1e-07 AD=1.4e-14 AS=1.15e-14 PD=4.8e-07 PS=4.3e-07 $X=127300 $Y=57665 $D=1
M498 GND 384 390 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.4e-14 AS=1.4e-14 PD=4.8e-07 PS=4.8e-07 $X=127680 $Y=54585 $D=1
M499 GND 384 392 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.4e-14 AS=1.4e-14 PD=4.8e-07 PS=4.8e-07 $X=127680 $Y=57665 $D=1
M500 GND RESET 193 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.2e-14 AS=1.2e-14 PD=4.4e-07 PS=4.4e-07 $X=127905 $Y=49225 $D=1
M501 390 165 GND GND NMOS_VTL L=5e-08 W=1e-07 AD=1.15e-14 AS=1.4e-14 PD=4.3e-07 PS=4.8e-07 $X=128060 $Y=54585 $D=1
M502 392 166 GND GND NMOS_VTL L=5e-08 W=1e-07 AD=1.15e-14 AS=1.4e-14 PD=4.3e-07 PS=4.8e-07 $X=128060 $Y=57665 $D=1
M503 GND 191 192 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.2e-14 AS=1.2e-14 PD=4.4e-07 PS=4.4e-07 $X=128765 $Y=49225 $D=1
M504 394 194 390 GND NMOS_VTL L=5e-08 W=9e-08 AD=1.08e-14 AS=1.125e-14 PD=4.2e-07 PS=4.3e-07 $X=128800 $Y=54585 $D=1
M505 395 195 392 GND NMOS_VTL L=5e-08 W=9e-08 AD=1.08e-14 AS=1.125e-14 PD=4.2e-07 PS=4.3e-07 $X=128800 $Y=57665 $D=1
M506 617 165 394 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.4e-14 AS=1.15e-14 PD=4.8e-07 PS=4.3e-07 $X=129530 $Y=54585 $D=1
M507 618 166 395 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.4e-14 AS=1.15e-14 PD=4.8e-07 PS=4.3e-07 $X=129530 $Y=57665 $D=1
M508 GND CLK_MAIN 191 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.2e-14 AS=1.2e-14 PD=4.4e-07 PS=4.4e-07 $X=129625 $Y=49225 $D=1
M509 619 381 617 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.4e-14 AS=1.4e-14 PD=4.8e-07 PS=4.8e-07 $X=129910 $Y=54585 $D=1
M510 620 381 618 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.4e-14 AS=1.4e-14 PD=4.8e-07 PS=4.8e-07 $X=129910 $Y=57665 $D=1
M511 GND 201 384 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.2e-14 AS=1.2e-14 PD=4.4e-07 PS=4.4e-07 $X=130020 $Y=62980 $D=1
M512 GND 201 200 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.2e-14 AS=1.2e-14 PD=4.4e-07 PS=4.4e-07 $X=130020 $Y=63840 $D=1
M513 621 200 201 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.5e-14 AS=1.2e-14 PD=5e-07 PS=4.4e-07 $X=130020 $Y=64700 $D=1
M514 622 198 621 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.4e-14 AS=1.5e-14 PD=4.8e-07 PS=5e-07 $X=130020 $Y=65100 $D=1
M515 GND 197 622 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.2e-14 AS=1.4e-14 PD=4.4e-07 PS=4.8e-07 $X=130020 $Y=65480 $D=1
M516 GND RESET 198 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.2e-14 AS=1.2e-14 PD=4.4e-07 PS=4.4e-07 $X=130020 $Y=66360 $D=1
M517 GND 197 196 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.2e-14 AS=1.2e-14 PD=4.4e-07 PS=4.4e-07 $X=130020 $Y=67220 $D=1
M518 GND CLK_MAIN 197 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.2e-14 AS=1.2e-14 PD=4.4e-07 PS=4.4e-07 $X=130020 $Y=68080 $D=1
M519 202 196 201 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.2e-14 AS=1.2e-14 PD=4.4e-07 PS=4.4e-07 $X=130020 $Y=68940 $D=1
M520 623 196 GND GND NMOS_VTL L=5e-08 W=1e-07 AD=1.4e-14 AS=1.2e-14 PD=4.8e-07 PS=4.4e-07 $X=130020 $Y=69800 $D=1
M521 199 202 623 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.2e-14 AS=1.4e-14 PD=4.4e-07 PS=4.8e-07 $X=130020 $Y=70180 $D=1
M522 624 198 202 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.5e-14 AS=1.2e-14 PD=5e-07 PS=4.4e-07 $X=130020 $Y=71040 $D=1
M523 GND 199 624 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.2e-14 AS=1.5e-14 PD=4.4e-07 PS=5e-07 $X=130020 $Y=71440 $D=1
M524 396 197 199 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.2e-14 AS=1.2e-14 PD=4.4e-07 PS=4.4e-07 $X=130020 $Y=72300 $D=1
M525 GND 397 396 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.2e-14 AS=1.2e-14 PD=4.4e-07 PS=4.4e-07 $X=130020 $Y=73160 $D=1
M526 GND B6 397 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.2e-14 AS=1.2e-14 PD=4.4e-07 PS=4.4e-07 $X=130020 $Y=74020 $D=1
M527 GND 384 619 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.15e-14 AS=1.4e-14 PD=4.3e-07 PS=4.8e-07 $X=130290 $Y=54585 $D=1
M528 GND 384 620 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.15e-14 AS=1.4e-14 PD=4.3e-07 PS=4.8e-07 $X=130290 $Y=57665 $D=1
M529 203 192 182 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.2e-14 AS=1.2e-14 PD=4.4e-07 PS=4.4e-07 $X=130485 $Y=49225 $D=1
M530 625 192 GND GND NMOS_VTL L=5e-08 W=1e-07 AD=1.4e-14 AS=1.2e-14 PD=4.8e-07 PS=4.4e-07 $X=131345 $Y=49225 $D=1
M531 208 394 GND GND NMOS_VTL L=5e-08 W=1e-07 AD=1.2e-14 AS=1.2e-14 PD=4.4e-07 PS=4.4e-07 $X=131395 $Y=55135 $D=1
M532 399 121 GND GND NMOS_VTL L=5e-08 W=1e-07 AD=1.35e-14 AS=1.15e-14 PD=4.7e-07 PS=4.3e-07 $X=131420 $Y=57305 $D=1
M533 205 203 625 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.2e-14 AS=1.4e-14 PD=4.4e-07 PS=4.8e-07 $X=131725 $Y=49225 $D=1
M534 SC6 399 206 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.4e-14 AS=1.2e-14 PD=4.8e-07 PS=4.4e-07 $X=132190 $Y=57305 $D=1
M535 GND 395 206 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.2e-14 AS=1.2e-14 PD=4.4e-07 PS=4.4e-07 $X=132400 $Y=58455 $D=1
M536 208 121 SC6 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.15e-14 AS=1.4e-14 PD=4.3e-07 PS=4.8e-07 $X=132570 $Y=57305 $D=1
M537 626 193 203 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.5e-14 AS=1.2e-14 PD=5e-07 PS=4.4e-07 $X=132585 $Y=49225 $D=1
M538 GND 205 626 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.2e-14 AS=1.5e-14 PD=4.4e-07 PS=5e-07 $X=132985 $Y=49225 $D=1
M539 400 191 205 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.2e-14 AS=1.2e-14 PD=4.4e-07 PS=4.4e-07 $X=133845 $Y=49225 $D=1
M540 GND 401 400 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.2e-14 AS=1.2e-14 PD=4.4e-07 PS=4.4e-07 $X=134705 $Y=49225 $D=1
M541 GND SC6 401 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.2e-14 AS=1.2e-14 PD=4.4e-07 PS=4.4e-07 $X=135565 $Y=49225 $D=1
M542 GND 404 403 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.2e-14 AS=1.2e-14 PD=4.4e-07 PS=4.4e-07 $X=136225 $Y=61795 $D=1
M543 GND 214 404 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.2e-14 AS=1.2e-14 PD=4.4e-07 PS=4.4e-07 $X=136225 $Y=62980 $D=1
M544 GND 214 213 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.2e-14 AS=1.2e-14 PD=4.4e-07 PS=4.4e-07 $X=136225 $Y=63840 $D=1
M545 627 213 214 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.5e-14 AS=1.2e-14 PD=5e-07 PS=4.4e-07 $X=136225 $Y=64700 $D=1
M546 628 211 627 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.4e-14 AS=1.5e-14 PD=4.8e-07 PS=5e-07 $X=136225 $Y=65100 $D=1
M547 GND 210 628 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.2e-14 AS=1.4e-14 PD=4.4e-07 PS=4.8e-07 $X=136225 $Y=65480 $D=1
M548 GND RESET 211 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.2e-14 AS=1.2e-14 PD=4.4e-07 PS=4.4e-07 $X=136225 $Y=66360 $D=1
M549 GND 210 209 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.2e-14 AS=1.2e-14 PD=4.4e-07 PS=4.4e-07 $X=136225 $Y=67220 $D=1
M550 GND CLK_MAIN 210 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.2e-14 AS=1.2e-14 PD=4.4e-07 PS=4.4e-07 $X=136225 $Y=68080 $D=1
M551 215 209 214 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.2e-14 AS=1.2e-14 PD=4.4e-07 PS=4.4e-07 $X=136225 $Y=68940 $D=1
M552 629 209 GND GND NMOS_VTL L=5e-08 W=1e-07 AD=1.4e-14 AS=1.2e-14 PD=4.8e-07 PS=4.4e-07 $X=136225 $Y=69800 $D=1
M553 212 215 629 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.2e-14 AS=1.4e-14 PD=4.4e-07 PS=4.8e-07 $X=136225 $Y=70180 $D=1
M554 630 211 215 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.5e-14 AS=1.2e-14 PD=5e-07 PS=4.4e-07 $X=136225 $Y=71040 $D=1
M555 GND 212 630 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.2e-14 AS=1.5e-14 PD=4.4e-07 PS=5e-07 $X=136225 $Y=71440 $D=1
M556 405 210 212 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.2e-14 AS=1.2e-14 PD=4.4e-07 PS=4.4e-07 $X=136225 $Y=72300 $D=1
M557 GND 406 405 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.2e-14 AS=1.2e-14 PD=4.4e-07 PS=4.4e-07 $X=136225 $Y=73160 $D=1
M558 GND A7 406 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.2e-14 AS=1.2e-14 PD=4.4e-07 PS=4.4e-07 $X=136225 $Y=74020 $D=1
M559 GND 403 408 GND NMOS_VTL L=5e-08 W=1.15e-07 AD=1.61e-14 AS=1.3225e-14 PD=5.1e-07 PS=4.6e-07 $X=136860 $Y=54555 $D=1
M560 GND 403 410 GND NMOS_VTL L=5e-08 W=1.15e-07 AD=1.61e-14 AS=1.3225e-14 PD=5.1e-07 PS=4.6e-07 $X=136860 $Y=57635 $D=1
M561 GND 216 S7 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.2e-14 AS=1.2e-14 PD=4.4e-07 PS=4.4e-07 $X=136905 $Y=49225 $D=1
M562 408 407 GND GND NMOS_VTL L=5e-08 W=1.15e-07 AD=1.61e-14 AS=1.61e-14 PD=5.1e-07 PS=5.1e-07 $X=137240 $Y=54555 $D=1
M563 410 407 GND GND NMOS_VTL L=5e-08 W=1.15e-07 AD=1.61e-14 AS=1.61e-14 PD=5.1e-07 PS=5.1e-07 $X=137240 $Y=57635 $D=1
M564 223 194 408 GND NMOS_VTL L=5e-08 W=1.15e-07 AD=1.61e-14 AS=1.61e-14 PD=5.1e-07 PS=5.1e-07 $X=137620 $Y=54555 $D=1
M565 224 195 410 GND NMOS_VTL L=5e-08 W=1.15e-07 AD=1.61e-14 AS=1.61e-14 PD=5.1e-07 PS=5.1e-07 $X=137620 $Y=57635 $D=1
M566 GND 216 218 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.2e-14 AS=1.2e-14 PD=4.4e-07 PS=4.4e-07 $X=137765 $Y=49225 $D=1
M567 631 403 223 GND NMOS_VTL L=5e-08 W=1.15e-07 AD=1.61e-14 AS=1.61e-14 PD=5.1e-07 PS=5.1e-07 $X=138000 $Y=54555 $D=1
M568 632 403 224 GND NMOS_VTL L=5e-08 W=1.15e-07 AD=1.61e-14 AS=1.61e-14 PD=5.1e-07 PS=5.1e-07 $X=138000 $Y=57635 $D=1
M569 GND 407 631 GND NMOS_VTL L=5e-08 W=1.15e-07 AD=1.3225e-14 AS=1.61e-14 PD=4.6e-07 PS=5.1e-07 $X=138380 $Y=54555 $D=1
M570 GND 407 632 GND NMOS_VTL L=5e-08 W=1.15e-07 AD=1.3225e-14 AS=1.61e-14 PD=4.6e-07 PS=5.1e-07 $X=138380 $Y=57635 $D=1
M571 633 218 216 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.5e-14 AS=1.2e-14 PD=5e-07 PS=4.4e-07 $X=138625 $Y=49225 $D=1
M572 634 222 633 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.4e-14 AS=1.5e-14 PD=4.8e-07 PS=5e-07 $X=139025 $Y=49225 $D=1
M573 413 403 GND GND NMOS_VTL L=5e-08 W=1e-07 AD=1.4e-14 AS=1.15e-14 PD=4.8e-07 PS=4.3e-07 $X=139100 $Y=54585 $D=1
M574 415 403 GND GND NMOS_VTL L=5e-08 W=1e-07 AD=1.4e-14 AS=1.15e-14 PD=4.8e-07 PS=4.3e-07 $X=139100 $Y=57665 $D=1
M575 GND 220 634 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.2e-14 AS=1.4e-14 PD=4.4e-07 PS=4.8e-07 $X=139405 $Y=49225 $D=1
M576 GND 407 413 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.4e-14 AS=1.4e-14 PD=4.8e-07 PS=4.8e-07 $X=139480 $Y=54585 $D=1
M577 GND 407 415 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.4e-14 AS=1.4e-14 PD=4.8e-07 PS=4.8e-07 $X=139480 $Y=57665 $D=1
M578 413 194 GND GND NMOS_VTL L=5e-08 W=1e-07 AD=1.15e-14 AS=1.4e-14 PD=4.3e-07 PS=4.8e-07 $X=139860 $Y=54585 $D=1
M579 415 195 GND GND NMOS_VTL L=5e-08 W=1e-07 AD=1.15e-14 AS=1.4e-14 PD=4.3e-07 PS=4.8e-07 $X=139860 $Y=57665 $D=1
M580 GND RESET 222 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.2e-14 AS=1.2e-14 PD=4.4e-07 PS=4.4e-07 $X=140285 $Y=49225 $D=1
M581 237 223 413 GND NMOS_VTL L=5e-08 W=9e-08 AD=1.08e-14 AS=1.125e-14 PD=4.2e-07 PS=4.3e-07 $X=140600 $Y=54585 $D=1
M582 234 224 415 GND NMOS_VTL L=5e-08 W=9e-08 AD=1.08e-14 AS=1.125e-14 PD=4.2e-07 PS=4.3e-07 $X=140600 $Y=57665 $D=1
M583 GND 220 221 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.2e-14 AS=1.2e-14 PD=4.4e-07 PS=4.4e-07 $X=141145 $Y=49225 $D=1
M584 635 194 237 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.4e-14 AS=1.15e-14 PD=4.8e-07 PS=4.3e-07 $X=141330 $Y=54585 $D=1
M585 636 195 234 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.4e-14 AS=1.15e-14 PD=4.8e-07 PS=4.3e-07 $X=141330 $Y=57665 $D=1
M586 641 403 635 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.4e-14 AS=1.4e-14 PD=4.8e-07 PS=4.8e-07 $X=141710 $Y=54585 $D=1
M587 642 403 636 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.4e-14 AS=1.4e-14 PD=4.8e-07 PS=4.8e-07 $X=141710 $Y=57665 $D=1
M588 GND 417 407 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.2e-14 AS=1.2e-14 PD=4.4e-07 PS=4.4e-07 $X=141745 $Y=61795 $D=1
M589 GND 230 417 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.2e-14 AS=1.2e-14 PD=4.4e-07 PS=4.4e-07 $X=141745 $Y=62980 $D=1
M590 GND 230 229 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.2e-14 AS=1.2e-14 PD=4.4e-07 PS=4.4e-07 $X=141745 $Y=63840 $D=1
M591 637 229 230 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.5e-14 AS=1.2e-14 PD=5e-07 PS=4.4e-07 $X=141745 $Y=64700 $D=1
M592 638 227 637 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.4e-14 AS=1.5e-14 PD=4.8e-07 PS=5e-07 $X=141745 $Y=65100 $D=1
M593 GND 226 638 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.2e-14 AS=1.4e-14 PD=4.4e-07 PS=4.8e-07 $X=141745 $Y=65480 $D=1
M594 GND RESET 227 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.2e-14 AS=1.2e-14 PD=4.4e-07 PS=4.4e-07 $X=141745 $Y=66360 $D=1
M595 GND 226 225 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.2e-14 AS=1.2e-14 PD=4.4e-07 PS=4.4e-07 $X=141745 $Y=67220 $D=1
M596 GND CLK_MAIN 226 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.2e-14 AS=1.2e-14 PD=4.4e-07 PS=4.4e-07 $X=141745 $Y=68080 $D=1
M597 231 225 230 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.2e-14 AS=1.2e-14 PD=4.4e-07 PS=4.4e-07 $X=141745 $Y=68940 $D=1
M598 639 225 GND GND NMOS_VTL L=5e-08 W=1e-07 AD=1.4e-14 AS=1.2e-14 PD=4.8e-07 PS=4.4e-07 $X=141745 $Y=69800 $D=1
M599 228 231 639 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.2e-14 AS=1.4e-14 PD=4.4e-07 PS=4.8e-07 $X=141745 $Y=70180 $D=1
M600 640 227 231 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.5e-14 AS=1.2e-14 PD=5e-07 PS=4.4e-07 $X=141745 $Y=71040 $D=1
M601 GND 228 640 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.2e-14 AS=1.5e-14 PD=4.4e-07 PS=5e-07 $X=141745 $Y=71440 $D=1
M602 418 226 228 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.2e-14 AS=1.2e-14 PD=4.4e-07 PS=4.4e-07 $X=141745 $Y=72300 $D=1
M603 GND 419 418 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.2e-14 AS=1.2e-14 PD=4.4e-07 PS=4.4e-07 $X=141745 $Y=73160 $D=1
M604 GND B7 419 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.2e-14 AS=1.2e-14 PD=4.4e-07 PS=4.4e-07 $X=141745 $Y=74020 $D=1
M605 GND CLK_MAIN 220 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.2e-14 AS=1.2e-14 PD=4.4e-07 PS=4.4e-07 $X=142005 $Y=49225 $D=1
M606 GND 407 641 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.15e-14 AS=1.4e-14 PD=4.3e-07 PS=4.8e-07 $X=142090 $Y=54585 $D=1
M607 GND 407 642 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.15e-14 AS=1.4e-14 PD=4.3e-07 PS=4.8e-07 $X=142090 $Y=57665 $D=1
M608 233 221 216 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.2e-14 AS=1.2e-14 PD=4.4e-07 PS=4.4e-07 $X=142865 $Y=49225 $D=1
M609 421 121 GND GND NMOS_VTL L=5e-08 W=1e-07 AD=1.35e-14 AS=1.15e-14 PD=4.7e-07 PS=4.3e-07 $X=143220 $Y=57305 $D=1
M610 643 221 GND GND NMOS_VTL L=5e-08 W=1e-07 AD=1.4e-14 AS=1.2e-14 PD=4.8e-07 PS=4.4e-07 $X=143725 $Y=49225 $D=1
M611 SC7 421 234 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.4e-14 AS=1.2e-14 PD=4.8e-07 PS=4.4e-07 $X=143990 $Y=57305 $D=1
M612 236 233 643 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.2e-14 AS=1.4e-14 PD=4.4e-07 PS=4.8e-07 $X=144105 $Y=49225 $D=1
M613 237 121 SC7 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.15e-14 AS=1.4e-14 PD=4.3e-07 PS=4.8e-07 $X=144370 $Y=57305 $D=1
M614 644 222 233 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.5e-14 AS=1.2e-14 PD=5e-07 PS=4.4e-07 $X=144965 $Y=49225 $D=1
M615 GND 236 644 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.2e-14 AS=1.5e-14 PD=4.4e-07 PS=5e-07 $X=145365 $Y=49225 $D=1
M616 423 220 236 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.2e-14 AS=1.2e-14 PD=4.4e-07 PS=4.4e-07 $X=146225 $Y=49225 $D=1
M617 422 121 GND GND NMOS_VTL L=5e-08 W=1e-07 AD=1.35e-14 AS=1.15e-14 PD=4.7e-07 PS=4.3e-07 $X=146325 $Y=57280 $D=1
M618 GND 424 423 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.2e-14 AS=1.2e-14 PD=4.4e-07 PS=4.4e-07 $X=147085 $Y=49225 $D=1
M619 C7_OUT 422 224 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.4e-14 AS=1.2e-14 PD=4.8e-07 PS=4.4e-07 $X=147095 $Y=57280 $D=1
M620 223 121 C7_OUT GND NMOS_VTL L=5e-08 W=1e-07 AD=1.15e-14 AS=1.4e-14 PD=4.3e-07 PS=4.8e-07 $X=147475 $Y=57280 $D=1
M621 GND SC7 424 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.2e-14 AS=1.2e-14 PD=4.4e-07 PS=4.4e-07 $X=147945 $Y=49225 $D=1
M622 426 C7_OUT GND GND NMOS_VTL L=5e-08 W=1e-07 AD=1.2e-14 AS=1.2e-14 PD=4.4e-07 PS=4.4e-07 $X=150115 $Y=57685 $D=1
M623 427 426 GND GND NMOS_VTL L=5e-08 W=1e-07 AD=1.2e-14 AS=1.2e-14 PD=4.4e-07 PS=4.4e-07 $X=150115 $Y=58545 $D=1
M624 245 243 427 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.2e-14 AS=1.2e-14 PD=4.4e-07 PS=4.4e-07 $X=150115 $Y=59405 $D=1
M625 645 245 GND GND NMOS_VTL L=5e-08 W=1e-07 AD=1.5e-14 AS=1.2e-14 PD=5e-07 PS=4.4e-07 $X=150115 $Y=60265 $D=1
M626 246 242 645 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.2e-14 AS=1.5e-14 PD=4.4e-07 PS=5e-07 $X=150115 $Y=60665 $D=1
M627 646 246 245 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.4e-14 AS=1.2e-14 PD=4.8e-07 PS=4.4e-07 $X=150115 $Y=61525 $D=1
M628 GND 239 646 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.2e-14 AS=1.4e-14 PD=4.4e-07 PS=4.8e-07 $X=150115 $Y=61905 $D=1
M629 241 239 246 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.2e-14 AS=1.2e-14 PD=4.4e-07 PS=4.4e-07 $X=150115 $Y=62765 $D=1
M630 243 CLK_MAIN GND GND NMOS_VTL L=5e-08 W=1e-07 AD=1.2e-14 AS=1.2e-14 PD=4.4e-07 PS=4.4e-07 $X=150115 $Y=63625 $D=1
M631 239 243 GND GND NMOS_VTL L=5e-08 W=1e-07 AD=1.2e-14 AS=1.2e-14 PD=4.4e-07 PS=4.4e-07 $X=150115 $Y=64485 $D=1
M632 242 RESET GND GND NMOS_VTL L=5e-08 W=1e-07 AD=1.2e-14 AS=1.2e-14 PD=4.4e-07 PS=4.4e-07 $X=150115 $Y=65345 $D=1
M633 647 243 GND GND NMOS_VTL L=5e-08 W=1e-07 AD=1.4e-14 AS=1.2e-14 PD=4.8e-07 PS=4.4e-07 $X=150115 $Y=66225 $D=1
M634 648 242 647 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.5e-14 AS=1.4e-14 PD=5e-07 PS=4.8e-07 $X=150115 $Y=66605 $D=1
M635 241 240 648 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.2e-14 AS=1.5e-14 PD=4.4e-07 PS=5e-07 $X=150115 $Y=67005 $D=1
M636 240 241 GND GND NMOS_VTL L=5e-08 W=1e-07 AD=1.2e-14 AS=1.2e-14 PD=4.4e-07 PS=4.4e-07 $X=150115 $Y=67865 $D=1
M637 Cout 241 GND GND NMOS_VTL L=5e-08 W=1e-07 AD=1.2e-14 AS=1.2e-14 PD=4.4e-07 PS=4.4e-07 $X=150115 $Y=68725 $D=1
M638 VDD 5 S0 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 $X=49850 $Y=50125 $D=0
M639 VDD 5 6 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 $X=50710 $Y=50125 $D=0
M640 VDD 248 253 VDD PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=2.07e-14 PD=6.4e-07 PS=5.9e-07 $X=50990 $Y=55935 $D=0
M641 VDD 248 255 VDD PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=2.07e-14 PD=6.4e-07 PS=5.9e-07 $X=50990 $Y=58855 $D=0
M642 VDD 10 248 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 $X=51350 $Y=62980 $D=0
M643 VDD 10 9 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 $X=51350 $Y=63840 $D=0
M644 10 9 13 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=2.4e-14 AS=1.92e-14 PD=6.2e-07 PS=5.6e-07 $X=51350 $Y=64700 $D=0
M645 13 7 10 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=2.4e-14 AS=2.4e-14 PD=6.2e-07 PS=6.2e-07 $X=51350 $Y=65100 $D=0
M646 VDD 3 13 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=1.92e-14 AS=2.4e-14 PD=5.6e-07 PS=6.2e-07 $X=51350 $Y=65500 $D=0
M647 VDD RESET 7 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 $X=51350 $Y=66360 $D=0
M648 VDD 4 3 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 $X=51350 $Y=67220 $D=0
M649 VDD CLK_MAIN 4 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 $X=51350 $Y=68080 $D=0
M650 11 4 10 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 $X=51350 $Y=68940 $D=0
M651 428 4 VDD VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=2.24e-14 AS=1.92e-14 PD=6e-07 PS=5.6e-07 $X=51350 $Y=69800 $D=0
M652 8 11 428 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=1.92e-14 AS=2.24e-14 PD=5.6e-07 PS=6e-07 $X=51350 $Y=70180 $D=0
M653 11 7 VDD VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=2.4e-14 AS=1.92e-14 PD=6.2e-07 PS=5.6e-07 $X=51350 $Y=71040 $D=0
M654 VDD 8 11 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=1.92e-14 AS=2.4e-14 PD=5.6e-07 PS=6.2e-07 $X=51350 $Y=71440 $D=0
M655 249 3 8 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 $X=51350 $Y=72300 $D=0
M656 VDD 250 249 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 $X=51350 $Y=73160 $D=0
M657 VDD A0 250 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 $X=51350 $Y=74020 $D=0
M658 253 251 VDD VDD PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=2.52e-14 PD=6.4e-07 PS=6.4e-07 $X=51370 $Y=55935 $D=0
M659 255 251 VDD VDD PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=2.52e-14 PD=6.4e-07 PS=6.4e-07 $X=51370 $Y=58855 $D=0
M660 5 6 12 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=2.4e-14 AS=1.92e-14 PD=6.2e-07 PS=5.6e-07 $X=51570 $Y=50125 $D=0
M661 19 VDD 253 VDD PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=2.52e-14 PD=6.4e-07 PS=6.4e-07 $X=51750 $Y=55935 $D=0
M662 20 GND 255 VDD PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=2.52e-14 PD=6.4e-07 PS=6.4e-07 $X=51750 $Y=58855 $D=0
M663 12 17 5 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=2.4e-14 AS=2.4e-14 PD=6.2e-07 PS=6.2e-07 $X=51970 $Y=50125 $D=0
M664 429 248 19 VDD PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=2.52e-14 PD=6.4e-07 PS=6.4e-07 $X=52130 $Y=55935 $D=0
M665 430 248 20 VDD PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=2.52e-14 PD=6.4e-07 PS=6.4e-07 $X=52130 $Y=58855 $D=0
M666 VDD 15 12 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=1.92e-14 AS=2.4e-14 PD=5.6e-07 PS=6.2e-07 $X=52370 $Y=50125 $D=0
M667 VDD 251 429 VDD PMOS_VTL L=5e-08 W=1.8e-07 AD=2.07e-14 AS=2.52e-14 PD=5.9e-07 PS=6.4e-07 $X=52510 $Y=55935 $D=0
M668 VDD 251 430 VDD PMOS_VTL L=5e-08 W=1.8e-07 AD=2.07e-14 AS=2.52e-14 PD=5.9e-07 PS=6.4e-07 $X=52510 $Y=58855 $D=0
M669 VDD RESET 17 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 $X=53230 $Y=50125 $D=0
M670 258 248 VDD VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=2.24e-14 AS=1.84e-14 PD=6e-07 PS=5.5e-07 $X=53230 $Y=55935 $D=0
M671 260 248 VDD VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=2.24e-14 AS=1.84e-14 PD=6e-07 PS=5.5e-07 $X=53230 $Y=58855 $D=0
M672 VDD 251 258 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=2.24e-14 AS=2.24e-14 PD=6e-07 PS=6e-07 $X=53610 $Y=55935 $D=0
M673 VDD 251 260 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=2.24e-14 AS=2.24e-14 PD=6e-07 PS=6e-07 $X=53610 $Y=58855 $D=0
M674 258 VDD VDD VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=1.84e-14 AS=2.24e-14 PD=5.5e-07 PS=6e-07 $X=53990 $Y=55935 $D=0
M675 260 GND VDD VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=1.84e-14 AS=2.24e-14 PD=5.5e-07 PS=6e-07 $X=53990 $Y=58855 $D=0
M676 VDD 14 15 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 $X=54090 $Y=50125 $D=0
M677 261 19 258 VDD PMOS_VTL L=5e-08 W=1.4e-07 AD=1.68e-14 AS=1.75e-14 PD=5.2e-07 PS=5.3e-07 $X=54730 $Y=55935 $D=0
M678 262 20 260 VDD PMOS_VTL L=5e-08 W=1.4e-07 AD=1.68e-14 AS=1.75e-14 PD=5.2e-07 PS=5.3e-07 $X=54730 $Y=58855 $D=0
M679 VDD CLK_MAIN 14 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 $X=54950 $Y=50125 $D=0
M680 431 VDD 261 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=2.24e-14 AS=1.84e-14 PD=6e-07 PS=5.5e-07 $X=55460 $Y=55935 $D=0
M681 432 GND 262 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=2.24e-14 AS=1.84e-14 PD=6e-07 PS=5.5e-07 $X=55460 $Y=58855 $D=0
M682 23 14 5 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 $X=55810 $Y=50125 $D=0
M683 433 248 431 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=2.24e-14 AS=2.24e-14 PD=6e-07 PS=6e-07 $X=55840 $Y=55935 $D=0
M684 434 248 432 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=2.24e-14 AS=2.24e-14 PD=6e-07 PS=6e-07 $X=55840 $Y=58855 $D=0
M685 VDD 251 433 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=1.84e-14 AS=2.24e-14 PD=5.5e-07 PS=6e-07 $X=56220 $Y=55935 $D=0
M686 VDD 251 434 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=1.84e-14 AS=2.24e-14 PD=5.5e-07 PS=6e-07 $X=56220 $Y=58855 $D=0
M687 435 14 VDD VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=2.24e-14 AS=1.92e-14 PD=6e-07 PS=5.6e-07 $X=56670 $Y=50125 $D=0
M688 VDD 27 251 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 $X=56850 $Y=62980 $D=0
M689 VDD 27 26 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 $X=56850 $Y=63840 $D=0
M690 27 26 29 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=2.4e-14 AS=1.92e-14 PD=6.2e-07 PS=5.6e-07 $X=56850 $Y=64700 $D=0
M691 29 24 27 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=2.4e-14 AS=2.4e-14 PD=6.2e-07 PS=6.2e-07 $X=56850 $Y=65100 $D=0
M692 VDD 21 29 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=1.92e-14 AS=2.4e-14 PD=5.6e-07 PS=6.2e-07 $X=56850 $Y=65500 $D=0
M693 VDD RESET 24 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 $X=56850 $Y=66360 $D=0
M694 VDD 22 21 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 $X=56850 $Y=67220 $D=0
M695 VDD CLK_MAIN 22 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 $X=56850 $Y=68080 $D=0
M696 28 22 27 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 $X=56850 $Y=68940 $D=0
M697 436 22 VDD VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=2.24e-14 AS=1.92e-14 PD=6e-07 PS=5.6e-07 $X=56850 $Y=69800 $D=0
M698 25 28 436 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=1.92e-14 AS=2.24e-14 PD=5.6e-07 PS=6e-07 $X=56850 $Y=70180 $D=0
M699 28 24 VDD VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=2.4e-14 AS=1.92e-14 PD=6.2e-07 PS=5.6e-07 $X=56850 $Y=71040 $D=0
M700 VDD 25 28 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=1.92e-14 AS=2.4e-14 PD=5.6e-07 PS=6.2e-07 $X=56850 $Y=71440 $D=0
M701 263 21 25 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 $X=56850 $Y=72300 $D=0
M702 VDD 264 263 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 $X=56850 $Y=73160 $D=0
M703 VDD B0 264 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 $X=56850 $Y=74020 $D=0
M704 30 23 435 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=1.92e-14 AS=2.24e-14 PD=5.6e-07 PS=6e-07 $X=57050 $Y=50125 $D=0
M705 VDD 262 31 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 $X=57320 $Y=58455 $D=0
M706 266 GND VDD VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=1.84e-14 AS=1.84e-14 PD=5.5e-07 PS=5.5e-07 $X=57350 $Y=56315 $D=0
M707 23 17 VDD VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=2.4e-14 AS=1.92e-14 PD=6.2e-07 PS=5.6e-07 $X=57910 $Y=50125 $D=0
M708 SC0 GND 31 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=2.24e-14 AS=1.84e-14 PD=6e-07 PS=5.5e-07 $X=58120 $Y=56315 $D=0
M709 33 261 VDD VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 $X=58215 $Y=55295 $D=0
M710 VDD 30 23 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=1.92e-14 AS=2.4e-14 PD=5.6e-07 PS=6.2e-07 $X=58310 $Y=50125 $D=0
M711 33 266 SC0 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=1.84e-14 AS=2.24e-14 PD=5.5e-07 PS=6e-07 $X=58500 $Y=56315 $D=0
M712 267 15 30 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 $X=59170 $Y=50125 $D=0
M713 VDD 268 267 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 $X=60030 $Y=50125 $D=0
M714 VDD SC0 268 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 $X=60890 $Y=50125 $D=0
M715 VDD 36 S1 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 $X=62115 $Y=50125 $D=0
M716 VDD 270 276 VDD PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=2.07e-14 PD=6.4e-07 PS=5.9e-07 $X=62790 $Y=55935 $D=0
M717 VDD 270 278 VDD PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=2.07e-14 PD=6.4e-07 PS=5.9e-07 $X=62790 $Y=59015 $D=0
M718 VDD 36 39 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 $X=62975 $Y=50125 $D=0
M719 VDD 271 270 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 $X=63045 $Y=61790 $D=0
M720 VDD 41 271 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 $X=63055 $Y=62975 $D=0
M721 VDD 41 40 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 $X=63055 $Y=63835 $D=0
M722 41 40 43 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=2.4e-14 AS=1.92e-14 PD=6.2e-07 PS=5.6e-07 $X=63055 $Y=64695 $D=0
M723 43 37 41 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=2.4e-14 AS=2.4e-14 PD=6.2e-07 PS=6.2e-07 $X=63055 $Y=65095 $D=0
M724 VDD 34 43 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=1.92e-14 AS=2.4e-14 PD=5.6e-07 PS=6.2e-07 $X=63055 $Y=65495 $D=0
M725 VDD RESET 37 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 $X=63055 $Y=66355 $D=0
M726 VDD 35 34 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 $X=63055 $Y=67215 $D=0
M727 VDD CLK_MAIN 35 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 $X=63055 $Y=68075 $D=0
M728 42 35 41 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 $X=63055 $Y=68935 $D=0
M729 437 35 VDD VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=2.24e-14 AS=1.92e-14 PD=6e-07 PS=5.6e-07 $X=63055 $Y=69795 $D=0
M730 38 42 437 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=1.92e-14 AS=2.24e-14 PD=5.6e-07 PS=6e-07 $X=63055 $Y=70175 $D=0
M731 42 37 VDD VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=2.4e-14 AS=1.92e-14 PD=6.2e-07 PS=5.6e-07 $X=63055 $Y=71035 $D=0
M732 VDD 38 42 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=1.92e-14 AS=2.4e-14 PD=5.6e-07 PS=6.2e-07 $X=63055 $Y=71435 $D=0
M733 272 34 38 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 $X=63055 $Y=72295 $D=0
M734 VDD 273 272 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 $X=63055 $Y=73155 $D=0
M735 VDD A1 273 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 $X=63055 $Y=74015 $D=0
M736 276 274 VDD VDD PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=2.52e-14 PD=6.4e-07 PS=6.4e-07 $X=63170 $Y=55935 $D=0
M737 278 274 VDD VDD PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=2.52e-14 PD=6.4e-07 PS=6.4e-07 $X=63170 $Y=59015 $D=0
M738 48 19 276 VDD PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=2.52e-14 PD=6.4e-07 PS=6.4e-07 $X=63550 $Y=55935 $D=0
M739 49 20 278 VDD PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=2.52e-14 PD=6.4e-07 PS=6.4e-07 $X=63550 $Y=59015 $D=0
M740 36 39 44 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=2.4e-14 AS=1.92e-14 PD=6.2e-07 PS=5.6e-07 $X=63835 $Y=50125 $D=0
M741 438 270 48 VDD PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=2.52e-14 PD=6.4e-07 PS=6.4e-07 $X=63930 $Y=55935 $D=0
M742 439 270 49 VDD PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=2.52e-14 PD=6.4e-07 PS=6.4e-07 $X=63930 $Y=59015 $D=0
M743 44 47 36 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=2.4e-14 AS=2.4e-14 PD=6.2e-07 PS=6.2e-07 $X=64235 $Y=50125 $D=0
M744 VDD 274 438 VDD PMOS_VTL L=5e-08 W=1.8e-07 AD=2.07e-14 AS=2.52e-14 PD=5.9e-07 PS=6.4e-07 $X=64310 $Y=55935 $D=0
M745 VDD 274 439 VDD PMOS_VTL L=5e-08 W=1.8e-07 AD=2.07e-14 AS=2.52e-14 PD=5.9e-07 PS=6.4e-07 $X=64310 $Y=59015 $D=0
M746 VDD 46 44 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=1.92e-14 AS=2.4e-14 PD=5.6e-07 PS=6.2e-07 $X=64635 $Y=50125 $D=0
M747 281 270 VDD VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=2.24e-14 AS=1.84e-14 PD=6e-07 PS=5.5e-07 $X=65030 $Y=55935 $D=0
M748 283 270 VDD VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=2.24e-14 AS=1.84e-14 PD=6e-07 PS=5.5e-07 $X=65030 $Y=59015 $D=0
M749 VDD 274 281 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=2.24e-14 AS=2.24e-14 PD=6e-07 PS=6e-07 $X=65410 $Y=55935 $D=0
M750 VDD 274 283 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=2.24e-14 AS=2.24e-14 PD=6e-07 PS=6e-07 $X=65410 $Y=59015 $D=0
M751 VDD RESET 47 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 $X=65495 $Y=50125 $D=0
M752 281 19 VDD VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=1.84e-14 AS=2.24e-14 PD=5.5e-07 PS=6e-07 $X=65790 $Y=55935 $D=0
M753 283 20 VDD VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=1.84e-14 AS=2.24e-14 PD=5.5e-07 PS=6e-07 $X=65790 $Y=59015 $D=0
M754 VDD 45 46 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 $X=66355 $Y=50125 $D=0
M755 62 48 281 VDD PMOS_VTL L=5e-08 W=1.4e-07 AD=1.68e-14 AS=1.75e-14 PD=5.2e-07 PS=5.3e-07 $X=66530 $Y=55935 $D=0
M756 60 49 283 VDD PMOS_VTL L=5e-08 W=1.4e-07 AD=1.68e-14 AS=1.75e-14 PD=5.2e-07 PS=5.3e-07 $X=66530 $Y=59015 $D=0
M757 VDD CLK_MAIN 45 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 $X=67215 $Y=50125 $D=0
M758 440 19 62 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=2.24e-14 AS=1.84e-14 PD=6e-07 PS=5.5e-07 $X=67260 $Y=55935 $D=0
M759 441 20 60 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=2.24e-14 AS=1.84e-14 PD=6e-07 PS=5.5e-07 $X=67260 $Y=59015 $D=0
M760 442 270 440 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=2.24e-14 AS=2.24e-14 PD=6e-07 PS=6e-07 $X=67640 $Y=55935 $D=0
M761 443 270 441 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=2.24e-14 AS=2.24e-14 PD=6e-07 PS=6e-07 $X=67640 $Y=59015 $D=0
M762 VDD 274 442 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=1.84e-14 AS=2.24e-14 PD=5.5e-07 PS=6e-07 $X=68020 $Y=55935 $D=0
M763 VDD 274 443 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=1.84e-14 AS=2.24e-14 PD=5.5e-07 PS=6e-07 $X=68020 $Y=59015 $D=0
M764 57 45 36 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 $X=68075 $Y=50125 $D=0
M765 VDD 284 274 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 $X=68565 $Y=61790 $D=0
M766 VDD 55 284 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 $X=68575 $Y=62975 $D=0
M767 VDD 55 54 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 $X=68575 $Y=63835 $D=0
M768 55 54 58 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=2.4e-14 AS=1.92e-14 PD=6.2e-07 PS=5.6e-07 $X=68575 $Y=64695 $D=0
M769 58 52 55 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=2.4e-14 AS=2.4e-14 PD=6.2e-07 PS=6.2e-07 $X=68575 $Y=65095 $D=0
M770 VDD 50 58 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=1.92e-14 AS=2.4e-14 PD=5.6e-07 PS=6.2e-07 $X=68575 $Y=65495 $D=0
M771 VDD RESET 52 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 $X=68575 $Y=66355 $D=0
M772 VDD 51 50 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 $X=68575 $Y=67215 $D=0
M773 VDD CLK_MAIN 51 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 $X=68575 $Y=68075 $D=0
M774 56 51 55 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 $X=68575 $Y=68935 $D=0
M775 444 51 VDD VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=2.24e-14 AS=1.92e-14 PD=6e-07 PS=5.6e-07 $X=68575 $Y=69795 $D=0
M776 53 56 444 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=1.92e-14 AS=2.24e-14 PD=5.6e-07 PS=6e-07 $X=68575 $Y=70175 $D=0
M777 56 52 VDD VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=2.4e-14 AS=1.92e-14 PD=6.2e-07 PS=5.6e-07 $X=68575 $Y=71035 $D=0
M778 VDD 53 56 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=1.92e-14 AS=2.4e-14 PD=5.6e-07 PS=6.2e-07 $X=68575 $Y=71435 $D=0
M779 285 50 53 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 $X=68575 $Y=72295 $D=0
M780 VDD 286 285 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 $X=68575 $Y=73155 $D=0
M781 VDD B1 286 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 $X=68575 $Y=74015 $D=0
M782 445 45 VDD VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=2.24e-14 AS=1.92e-14 PD=6e-07 PS=5.6e-07 $X=68935 $Y=50125 $D=0
M783 288 GND VDD VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=1.84e-14 AS=1.84e-14 PD=5.5e-07 PS=5.5e-07 $X=69150 $Y=56475 $D=0
M784 59 57 445 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=1.92e-14 AS=2.24e-14 PD=5.6e-07 PS=6e-07 $X=69315 $Y=50125 $D=0
M785 SC1 GND 60 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=2.24e-14 AS=1.84e-14 PD=6e-07 PS=5.5e-07 $X=69920 $Y=56475 $D=0
M786 57 47 VDD VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=2.4e-14 AS=1.92e-14 PD=6.2e-07 PS=5.6e-07 $X=70175 $Y=50125 $D=0
M787 62 288 SC1 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=1.84e-14 AS=2.24e-14 PD=5.5e-07 PS=6e-07 $X=70300 $Y=56475 $D=0
M788 VDD 59 57 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=1.92e-14 AS=2.4e-14 PD=5.6e-07 PS=6.2e-07 $X=70575 $Y=50125 $D=0
M789 289 46 59 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 $X=71435 $Y=50125 $D=0
M790 VDD 290 289 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 $X=72295 $Y=50125 $D=0
M791 VDD SC1 290 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 $X=73155 $Y=50125 $D=0
M792 VDD 67 S2 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 $X=74310 $Y=50125 $D=0
M793 VDD 292 297 VDD PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=2.07e-14 PD=6.4e-07 PS=5.9e-07 $X=74590 $Y=55935 $D=0
M794 VDD 292 299 VDD PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=2.07e-14 PD=6.4e-07 PS=5.9e-07 $X=74590 $Y=59015 $D=0
M795 VDD 69 292 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 $X=74950 $Y=62980 $D=0
M796 VDD 69 68 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 $X=74950 $Y=63840 $D=0
M797 69 68 72 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=2.4e-14 AS=1.92e-14 PD=6.2e-07 PS=5.6e-07 $X=74950 $Y=64700 $D=0
M798 72 65 69 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=2.4e-14 AS=2.4e-14 PD=6.2e-07 PS=6.2e-07 $X=74950 $Y=65100 $D=0
M799 VDD 63 72 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=1.92e-14 AS=2.4e-14 PD=5.6e-07 PS=6.2e-07 $X=74950 $Y=65500 $D=0
M800 VDD RESET 65 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 $X=74950 $Y=66360 $D=0
M801 VDD 64 63 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 $X=74950 $Y=67220 $D=0
M802 VDD CLK_MAIN 64 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 $X=74950 $Y=68080 $D=0
M803 70 64 69 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 $X=74950 $Y=68940 $D=0
M804 446 64 VDD VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=2.24e-14 AS=1.92e-14 PD=6e-07 PS=5.6e-07 $X=74950 $Y=69800 $D=0
M805 66 70 446 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=1.92e-14 AS=2.24e-14 PD=5.6e-07 PS=6e-07 $X=74950 $Y=70180 $D=0
M806 70 65 VDD VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=2.4e-14 AS=1.92e-14 PD=6.2e-07 PS=5.6e-07 $X=74950 $Y=71040 $D=0
M807 VDD 66 70 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=1.92e-14 AS=2.4e-14 PD=5.6e-07 PS=6.2e-07 $X=74950 $Y=71440 $D=0
M808 293 63 66 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 $X=74950 $Y=72300 $D=0
M809 VDD 294 293 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 $X=74950 $Y=73160 $D=0
M810 VDD A2 294 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 $X=74950 $Y=74020 $D=0
M811 297 295 VDD VDD PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=2.52e-14 PD=6.4e-07 PS=6.4e-07 $X=74970 $Y=55935 $D=0
M812 299 295 VDD VDD PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=2.52e-14 PD=6.4e-07 PS=6.4e-07 $X=74970 $Y=59015 $D=0
M813 VDD 67 71 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 $X=75170 $Y=50125 $D=0
M814 77 48 297 VDD PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=2.52e-14 PD=6.4e-07 PS=6.4e-07 $X=75350 $Y=55935 $D=0
M815 78 49 299 VDD PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=2.52e-14 PD=6.4e-07 PS=6.4e-07 $X=75350 $Y=59015 $D=0
M816 447 292 77 VDD PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=2.52e-14 PD=6.4e-07 PS=6.4e-07 $X=75730 $Y=55935 $D=0
M817 448 292 78 VDD PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=2.52e-14 PD=6.4e-07 PS=6.4e-07 $X=75730 $Y=59015 $D=0
M818 67 71 73 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=2.4e-14 AS=1.92e-14 PD=6.2e-07 PS=5.6e-07 $X=76030 $Y=50125 $D=0
M819 VDD 295 447 VDD PMOS_VTL L=5e-08 W=1.8e-07 AD=2.07e-14 AS=2.52e-14 PD=5.9e-07 PS=6.4e-07 $X=76110 $Y=55935 $D=0
M820 VDD 295 448 VDD PMOS_VTL L=5e-08 W=1.8e-07 AD=2.07e-14 AS=2.52e-14 PD=5.9e-07 PS=6.4e-07 $X=76110 $Y=59015 $D=0
M821 73 76 67 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=2.4e-14 AS=2.4e-14 PD=6.2e-07 PS=6.2e-07 $X=76430 $Y=50125 $D=0
M822 VDD 75 73 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=1.92e-14 AS=2.4e-14 PD=5.6e-07 PS=6.2e-07 $X=76830 $Y=50125 $D=0
M823 302 292 VDD VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=2.24e-14 AS=1.84e-14 PD=6e-07 PS=5.5e-07 $X=76830 $Y=55935 $D=0
M824 304 292 VDD VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=2.24e-14 AS=1.84e-14 PD=6e-07 PS=5.5e-07 $X=76830 $Y=59015 $D=0
M825 VDD 295 302 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=2.24e-14 AS=2.24e-14 PD=6e-07 PS=6e-07 $X=77210 $Y=55935 $D=0
M826 VDD 295 304 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=2.24e-14 AS=2.24e-14 PD=6e-07 PS=6e-07 $X=77210 $Y=59015 $D=0
M827 302 48 VDD VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=1.84e-14 AS=2.24e-14 PD=5.5e-07 PS=6e-07 $X=77590 $Y=55935 $D=0
M828 304 49 VDD VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=1.84e-14 AS=2.24e-14 PD=5.5e-07 PS=6e-07 $X=77590 $Y=59015 $D=0
M829 VDD RESET 76 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 $X=77690 $Y=50125 $D=0
M830 305 77 302 VDD PMOS_VTL L=5e-08 W=1.4e-07 AD=1.68e-14 AS=1.75e-14 PD=5.2e-07 PS=5.3e-07 $X=78330 $Y=55935 $D=0
M831 306 78 304 VDD PMOS_VTL L=5e-08 W=1.4e-07 AD=1.68e-14 AS=1.75e-14 PD=5.2e-07 PS=5.3e-07 $X=78330 $Y=59015 $D=0
M832 VDD 74 75 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 $X=78550 $Y=50125 $D=0
M833 449 48 305 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=2.24e-14 AS=1.84e-14 PD=6e-07 PS=5.5e-07 $X=79060 $Y=55935 $D=0
M834 450 49 306 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=2.24e-14 AS=1.84e-14 PD=6e-07 PS=5.5e-07 $X=79060 $Y=59015 $D=0
M835 VDD CLK_MAIN 74 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 $X=79410 $Y=50125 $D=0
M836 451 292 449 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=2.24e-14 AS=2.24e-14 PD=6e-07 PS=6e-07 $X=79440 $Y=55935 $D=0
M837 452 292 450 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=2.24e-14 AS=2.24e-14 PD=6e-07 PS=6e-07 $X=79440 $Y=59015 $D=0
M838 VDD 295 451 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=1.84e-14 AS=2.24e-14 PD=5.5e-07 PS=6e-07 $X=79820 $Y=55935 $D=0
M839 VDD 295 452 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=1.84e-14 AS=2.24e-14 PD=5.5e-07 PS=6e-07 $X=79820 $Y=59015 $D=0
M840 86 74 67 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 $X=80270 $Y=50125 $D=0
M841 VDD 84 295 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 $X=80450 $Y=62980 $D=0
M842 VDD 84 83 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 $X=80450 $Y=63840 $D=0
M843 84 83 87 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=2.4e-14 AS=1.92e-14 PD=6.2e-07 PS=5.6e-07 $X=80450 $Y=64700 $D=0
M844 87 81 84 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=2.4e-14 AS=2.4e-14 PD=6.2e-07 PS=6.2e-07 $X=80450 $Y=65100 $D=0
M845 VDD 79 87 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=1.92e-14 AS=2.4e-14 PD=5.6e-07 PS=6.2e-07 $X=80450 $Y=65500 $D=0
M846 VDD RESET 81 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 $X=80450 $Y=66360 $D=0
M847 VDD 80 79 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 $X=80450 $Y=67220 $D=0
M848 VDD CLK_MAIN 80 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 $X=80450 $Y=68080 $D=0
M849 85 80 84 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 $X=80450 $Y=68940 $D=0
M850 453 80 VDD VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=2.24e-14 AS=1.92e-14 PD=6e-07 PS=5.6e-07 $X=80450 $Y=69800 $D=0
M851 82 85 453 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=1.92e-14 AS=2.24e-14 PD=5.6e-07 PS=6e-07 $X=80450 $Y=70180 $D=0
M852 85 81 VDD VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=2.4e-14 AS=1.92e-14 PD=6.2e-07 PS=5.6e-07 $X=80450 $Y=71040 $D=0
M853 VDD 82 85 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=1.92e-14 AS=2.4e-14 PD=5.6e-07 PS=6.2e-07 $X=80450 $Y=71440 $D=0
M854 307 79 82 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 $X=80450 $Y=72300 $D=0
M855 VDD 308 307 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 $X=80450 $Y=73160 $D=0
M856 VDD B2 308 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 $X=80450 $Y=74020 $D=0
M857 VDD 306 88 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 $X=80920 $Y=58615 $D=0
M858 310 GND VDD VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=1.84e-14 AS=1.84e-14 PD=5.5e-07 PS=5.5e-07 $X=80950 $Y=56475 $D=0
M859 454 74 VDD VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=2.24e-14 AS=1.92e-14 PD=6e-07 PS=5.6e-07 $X=81130 $Y=50125 $D=0
M860 89 86 454 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=1.92e-14 AS=2.24e-14 PD=5.6e-07 PS=6e-07 $X=81510 $Y=50125 $D=0
M861 SC2 GND 88 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=2.24e-14 AS=1.84e-14 PD=6e-07 PS=5.5e-07 $X=81720 $Y=56475 $D=0
M862 91 305 VDD VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 $X=81815 $Y=55295 $D=0
M863 91 310 SC2 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=1.84e-14 AS=2.24e-14 PD=5.5e-07 PS=6e-07 $X=82100 $Y=56475 $D=0
M864 86 76 VDD VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=2.4e-14 AS=1.92e-14 PD=6.2e-07 PS=5.6e-07 $X=82370 $Y=50125 $D=0
M865 VDD 89 86 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=1.92e-14 AS=2.4e-14 PD=5.6e-07 PS=6.2e-07 $X=82770 $Y=50125 $D=0
M866 311 75 89 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 $X=83630 $Y=50125 $D=0
M867 VDD 312 311 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 $X=84490 $Y=50125 $D=0
M868 VDD SC2 312 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 $X=85350 $Y=50125 $D=0
M869 VDD 313 320 VDD PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=2.07e-14 PD=6.4e-07 PS=5.9e-07 $X=86390 $Y=55775 $D=0
M870 VDD 313 322 VDD PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=2.07e-14 PD=6.4e-07 PS=5.9e-07 $X=86390 $Y=58855 $D=0
M871 VDD 99 S3 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 $X=86575 $Y=50125 $D=0
M872 VDD 315 313 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 $X=86645 $Y=61795 $D=0
M873 VDD 97 315 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 $X=86655 $Y=62980 $D=0
M874 VDD 97 96 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 $X=86655 $Y=63840 $D=0
M875 97 96 100 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=2.4e-14 AS=1.92e-14 PD=6.2e-07 PS=5.6e-07 $X=86655 $Y=64700 $D=0
M876 100 94 97 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=2.4e-14 AS=2.4e-14 PD=6.2e-07 PS=6.2e-07 $X=86655 $Y=65100 $D=0
M877 VDD 92 100 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=1.92e-14 AS=2.4e-14 PD=5.6e-07 PS=6.2e-07 $X=86655 $Y=65500 $D=0
M878 VDD RESET 94 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 $X=86655 $Y=66360 $D=0
M879 VDD 93 92 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 $X=86655 $Y=67220 $D=0
M880 VDD CLK_MAIN 93 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 $X=86655 $Y=68080 $D=0
M881 98 93 97 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 $X=86655 $Y=68940 $D=0
M882 455 93 VDD VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=2.24e-14 AS=1.92e-14 PD=6e-07 PS=5.6e-07 $X=86655 $Y=69800 $D=0
M883 95 98 455 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=1.92e-14 AS=2.24e-14 PD=5.6e-07 PS=6e-07 $X=86655 $Y=70180 $D=0
M884 98 94 VDD VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=2.4e-14 AS=1.92e-14 PD=6.2e-07 PS=5.6e-07 $X=86655 $Y=71040 $D=0
M885 VDD 95 98 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=1.92e-14 AS=2.4e-14 PD=5.6e-07 PS=6.2e-07 $X=86655 $Y=71440 $D=0
M886 316 92 95 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 $X=86655 $Y=72300 $D=0
M887 VDD 317 316 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 $X=86655 $Y=73160 $D=0
M888 VDD A3 317 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 $X=86655 $Y=74020 $D=0
M889 320 318 VDD VDD PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=2.52e-14 PD=6.4e-07 PS=6.4e-07 $X=86770 $Y=55775 $D=0
M890 322 318 VDD VDD PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=2.52e-14 PD=6.4e-07 PS=6.4e-07 $X=86770 $Y=58855 $D=0
M891 106 77 320 VDD PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=2.52e-14 PD=6.4e-07 PS=6.4e-07 $X=87150 $Y=55775 $D=0
M892 107 78 322 VDD PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=2.52e-14 PD=6.4e-07 PS=6.4e-07 $X=87150 $Y=58855 $D=0
M893 VDD 99 101 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 $X=87435 $Y=50125 $D=0
M894 456 313 106 VDD PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=2.52e-14 PD=6.4e-07 PS=6.4e-07 $X=87530 $Y=55775 $D=0
M895 457 313 107 VDD PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=2.52e-14 PD=6.4e-07 PS=6.4e-07 $X=87530 $Y=58855 $D=0
M896 VDD 318 456 VDD PMOS_VTL L=5e-08 W=1.8e-07 AD=2.07e-14 AS=2.52e-14 PD=5.9e-07 PS=6.4e-07 $X=87910 $Y=55775 $D=0
M897 VDD 318 457 VDD PMOS_VTL L=5e-08 W=1.8e-07 AD=2.07e-14 AS=2.52e-14 PD=5.9e-07 PS=6.4e-07 $X=87910 $Y=58855 $D=0
M898 99 101 102 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=2.4e-14 AS=1.92e-14 PD=6.2e-07 PS=5.6e-07 $X=88295 $Y=50125 $D=0
M899 325 313 VDD VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=2.24e-14 AS=1.84e-14 PD=6e-07 PS=5.5e-07 $X=88630 $Y=55775 $D=0
M900 327 313 VDD VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=2.24e-14 AS=1.84e-14 PD=6e-07 PS=5.5e-07 $X=88630 $Y=58855 $D=0
M901 102 105 99 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=2.4e-14 AS=2.4e-14 PD=6.2e-07 PS=6.2e-07 $X=88695 $Y=50125 $D=0
M902 VDD 318 325 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=2.24e-14 AS=2.24e-14 PD=6e-07 PS=6e-07 $X=89010 $Y=55775 $D=0
M903 VDD 318 327 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=2.24e-14 AS=2.24e-14 PD=6e-07 PS=6e-07 $X=89010 $Y=58855 $D=0
M904 VDD 104 102 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=1.92e-14 AS=2.4e-14 PD=5.6e-07 PS=6.2e-07 $X=89095 $Y=50125 $D=0
M905 325 77 VDD VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=1.84e-14 AS=2.24e-14 PD=5.5e-07 PS=6e-07 $X=89390 $Y=55775 $D=0
M906 327 78 VDD VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=1.84e-14 AS=2.24e-14 PD=5.5e-07 PS=6e-07 $X=89390 $Y=58855 $D=0
M907 VDD RESET 105 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 $X=89955 $Y=50125 $D=0
M908 120 106 325 VDD PMOS_VTL L=5e-08 W=1.4e-07 AD=1.68e-14 AS=1.75e-14 PD=5.2e-07 PS=5.3e-07 $X=90130 $Y=55775 $D=0
M909 117 107 327 VDD PMOS_VTL L=5e-08 W=1.4e-07 AD=1.68e-14 AS=1.75e-14 PD=5.2e-07 PS=5.3e-07 $X=90130 $Y=58855 $D=0
M910 VDD 103 104 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 $X=90815 $Y=50125 $D=0
M911 458 77 120 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=2.24e-14 AS=1.84e-14 PD=6e-07 PS=5.5e-07 $X=90860 $Y=55775 $D=0
M912 459 78 117 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=2.24e-14 AS=1.84e-14 PD=6e-07 PS=5.5e-07 $X=90860 $Y=58855 $D=0
M913 460 313 458 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=2.24e-14 AS=2.24e-14 PD=6e-07 PS=6e-07 $X=91240 $Y=55775 $D=0
M914 461 313 459 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=2.24e-14 AS=2.24e-14 PD=6e-07 PS=6e-07 $X=91240 $Y=58855 $D=0
M915 VDD 318 460 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=1.84e-14 AS=2.24e-14 PD=5.5e-07 PS=6e-07 $X=91620 $Y=55775 $D=0
M916 VDD 318 461 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=1.84e-14 AS=2.24e-14 PD=5.5e-07 PS=6e-07 $X=91620 $Y=58855 $D=0
M917 VDD CLK_MAIN 103 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 $X=91675 $Y=50125 $D=0
M918 VDD 328 318 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 $X=92165 $Y=61795 $D=0
M919 VDD 113 328 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 $X=92175 $Y=62980 $D=0
M920 VDD 113 112 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 $X=92175 $Y=63840 $D=0
M921 113 112 115 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=2.4e-14 AS=1.92e-14 PD=6.2e-07 PS=5.6e-07 $X=92175 $Y=64700 $D=0
M922 115 110 113 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=2.4e-14 AS=2.4e-14 PD=6.2e-07 PS=6.2e-07 $X=92175 $Y=65100 $D=0
M923 VDD 108 115 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=1.92e-14 AS=2.4e-14 PD=5.6e-07 PS=6.2e-07 $X=92175 $Y=65500 $D=0
M924 VDD RESET 110 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 $X=92175 $Y=66360 $D=0
M925 VDD 109 108 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 $X=92175 $Y=67220 $D=0
M926 VDD CLK_MAIN 109 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 $X=92175 $Y=68080 $D=0
M927 114 109 113 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 $X=92175 $Y=68940 $D=0
M928 462 109 VDD VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=2.24e-14 AS=1.92e-14 PD=6e-07 PS=5.6e-07 $X=92175 $Y=69800 $D=0
M929 111 114 462 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=1.92e-14 AS=2.24e-14 PD=5.6e-07 PS=6e-07 $X=92175 $Y=70180 $D=0
M930 114 110 VDD VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=2.4e-14 AS=1.92e-14 PD=6.2e-07 PS=5.6e-07 $X=92175 $Y=71040 $D=0
M931 VDD 111 114 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=1.92e-14 AS=2.4e-14 PD=5.6e-07 PS=6.2e-07 $X=92175 $Y=71440 $D=0
M932 329 108 111 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 $X=92175 $Y=72300 $D=0
M933 VDD 330 329 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 $X=92175 $Y=73160 $D=0
M934 VDD B3 330 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 $X=92175 $Y=74020 $D=0
M935 116 103 99 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 $X=92535 $Y=50125 $D=0
M936 332 GND VDD VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=1.84e-14 AS=1.84e-14 PD=5.5e-07 PS=5.5e-07 $X=92750 $Y=56315 $D=0
M937 463 103 VDD VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=2.24e-14 AS=1.92e-14 PD=6e-07 PS=5.6e-07 $X=93395 $Y=50125 $D=0
M938 SC3 GND 117 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=2.24e-14 AS=1.84e-14 PD=6e-07 PS=5.5e-07 $X=93520 $Y=56315 $D=0
M939 119 116 463 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=1.92e-14 AS=2.24e-14 PD=5.6e-07 PS=6e-07 $X=93775 $Y=50125 $D=0
M940 120 332 SC3 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=1.84e-14 AS=2.24e-14 PD=5.5e-07 PS=6e-07 $X=93900 $Y=56315 $D=0
M941 116 105 VDD VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=2.4e-14 AS=1.92e-14 PD=6.2e-07 PS=5.6e-07 $X=94635 $Y=50125 $D=0
M942 VDD 119 116 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=1.92e-14 AS=2.4e-14 PD=5.6e-07 PS=6.2e-07 $X=95035 $Y=50125 $D=0
M943 333 GND VDD VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=1.84e-14 AS=1.84e-14 PD=5.5e-07 PS=5.5e-07 $X=95855 $Y=56290 $D=0
M944 334 104 119 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 $X=95895 $Y=50125 $D=0
M945 121 GND 107 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=2.24e-14 AS=1.84e-14 PD=6e-07 PS=5.5e-07 $X=96625 $Y=56290 $D=0
M946 VDD 335 334 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 $X=96755 $Y=50125 $D=0
M947 106 333 121 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=1.84e-14 AS=2.24e-14 PD=5.5e-07 PS=6e-07 $X=97005 $Y=56290 $D=0
M948 VDD SC3 335 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 $X=97615 $Y=50125 $D=0
M949 VDD 122 S4 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 $X=99550 $Y=50125 $D=0
M950 VDD 122 123 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 $X=100410 $Y=50125 $D=0
M951 122 123 126 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=2.4e-14 AS=1.92e-14 PD=6.2e-07 PS=5.6e-07 $X=101270 $Y=50125 $D=0
M952 VDD 337 342 VDD PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=2.07e-14 PD=6.4e-07 PS=5.9e-07 $X=101460 $Y=55935 $D=0
M953 VDD 337 344 VDD PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=2.07e-14 PD=6.4e-07 PS=5.9e-07 $X=101460 $Y=58855 $D=0
M954 126 135 122 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=2.4e-14 AS=2.4e-14 PD=6.2e-07 PS=6.2e-07 $X=101670 $Y=50125 $D=0
M955 VDD 130 337 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 $X=101820 $Y=62980 $D=0
M956 VDD 130 129 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 $X=101820 $Y=63840 $D=0
M957 130 129 132 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=2.4e-14 AS=1.92e-14 PD=6.2e-07 PS=5.6e-07 $X=101820 $Y=64700 $D=0
M958 132 127 130 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=2.4e-14 AS=2.4e-14 PD=6.2e-07 PS=6.2e-07 $X=101820 $Y=65100 $D=0
M959 VDD 124 132 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=1.92e-14 AS=2.4e-14 PD=5.6e-07 PS=6.2e-07 $X=101820 $Y=65500 $D=0
M960 VDD RESET 127 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 $X=101820 $Y=66360 $D=0
M961 VDD 125 124 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 $X=101820 $Y=67220 $D=0
M962 VDD CLK_MAIN 125 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 $X=101820 $Y=68080 $D=0
M963 131 125 130 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 $X=101820 $Y=68940 $D=0
M964 464 125 VDD VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=2.24e-14 AS=1.92e-14 PD=6e-07 PS=5.6e-07 $X=101820 $Y=69800 $D=0
M965 128 131 464 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=1.92e-14 AS=2.24e-14 PD=5.6e-07 PS=6e-07 $X=101820 $Y=70180 $D=0
M966 131 127 VDD VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=2.4e-14 AS=1.92e-14 PD=6.2e-07 PS=5.6e-07 $X=101820 $Y=71040 $D=0
M967 VDD 128 131 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=1.92e-14 AS=2.4e-14 PD=5.6e-07 PS=6.2e-07 $X=101820 $Y=71440 $D=0
M968 338 124 128 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 $X=101820 $Y=72300 $D=0
M969 VDD 339 338 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 $X=101820 $Y=73160 $D=0
M970 VDD A4 339 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 $X=101820 $Y=74020 $D=0
M971 342 340 VDD VDD PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=2.52e-14 PD=6.4e-07 PS=6.4e-07 $X=101840 $Y=55935 $D=0
M972 344 340 VDD VDD PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=2.52e-14 PD=6.4e-07 PS=6.4e-07 $X=101840 $Y=58855 $D=0
M973 VDD 134 126 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=1.92e-14 AS=2.4e-14 PD=5.6e-07 PS=6.2e-07 $X=102070 $Y=50125 $D=0
M974 136 VDD 342 VDD PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=2.52e-14 PD=6.4e-07 PS=6.4e-07 $X=102220 $Y=55935 $D=0
M975 137 GND 344 VDD PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=2.52e-14 PD=6.4e-07 PS=6.4e-07 $X=102220 $Y=58855 $D=0
M976 465 337 136 VDD PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=2.52e-14 PD=6.4e-07 PS=6.4e-07 $X=102600 $Y=55935 $D=0
M977 466 337 137 VDD PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=2.52e-14 PD=6.4e-07 PS=6.4e-07 $X=102600 $Y=58855 $D=0
M978 VDD RESET 135 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 $X=102930 $Y=50125 $D=0
M979 VDD 340 465 VDD PMOS_VTL L=5e-08 W=1.8e-07 AD=2.07e-14 AS=2.52e-14 PD=5.9e-07 PS=6.4e-07 $X=102980 $Y=55935 $D=0
M980 VDD 340 466 VDD PMOS_VTL L=5e-08 W=1.8e-07 AD=2.07e-14 AS=2.52e-14 PD=5.9e-07 PS=6.4e-07 $X=102980 $Y=58855 $D=0
M981 347 337 VDD VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=2.24e-14 AS=1.84e-14 PD=6e-07 PS=5.5e-07 $X=103700 $Y=55935 $D=0
M982 349 337 VDD VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=2.24e-14 AS=1.84e-14 PD=6e-07 PS=5.5e-07 $X=103700 $Y=58855 $D=0
M983 VDD 133 134 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 $X=103790 $Y=50125 $D=0
M984 VDD 340 347 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=2.24e-14 AS=2.24e-14 PD=6e-07 PS=6e-07 $X=104080 $Y=55935 $D=0
M985 VDD 340 349 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=2.24e-14 AS=2.24e-14 PD=6e-07 PS=6e-07 $X=104080 $Y=58855 $D=0
M986 347 VDD VDD VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=1.84e-14 AS=2.24e-14 PD=5.5e-07 PS=6e-07 $X=104460 $Y=55935 $D=0
M987 349 GND VDD VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=1.84e-14 AS=2.24e-14 PD=5.5e-07 PS=6e-07 $X=104460 $Y=58855 $D=0
M988 VDD CLK_MAIN 133 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 $X=104650 $Y=50125 $D=0
M989 350 136 347 VDD PMOS_VTL L=5e-08 W=1.4e-07 AD=1.68e-14 AS=1.75e-14 PD=5.2e-07 PS=5.3e-07 $X=105200 $Y=55935 $D=0
M990 351 137 349 VDD PMOS_VTL L=5e-08 W=1.4e-07 AD=1.68e-14 AS=1.75e-14 PD=5.2e-07 PS=5.3e-07 $X=105200 $Y=58855 $D=0
M991 139 133 122 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 $X=105510 $Y=50125 $D=0
M992 467 VDD 350 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=2.24e-14 AS=1.84e-14 PD=6e-07 PS=5.5e-07 $X=105930 $Y=55935 $D=0
M993 468 GND 351 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=2.24e-14 AS=1.84e-14 PD=6e-07 PS=5.5e-07 $X=105930 $Y=58855 $D=0
M994 469 337 467 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=2.24e-14 AS=2.24e-14 PD=6e-07 PS=6e-07 $X=106310 $Y=55935 $D=0
M995 470 337 468 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=2.24e-14 AS=2.24e-14 PD=6e-07 PS=6e-07 $X=106310 $Y=58855 $D=0
M996 471 133 VDD VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=2.24e-14 AS=1.92e-14 PD=6e-07 PS=5.6e-07 $X=106370 $Y=50125 $D=0
M997 VDD 340 469 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=1.84e-14 AS=2.24e-14 PD=5.5e-07 PS=6e-07 $X=106690 $Y=55935 $D=0
M998 VDD 340 470 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=1.84e-14 AS=2.24e-14 PD=5.5e-07 PS=6e-07 $X=106690 $Y=58855 $D=0
M999 146 139 471 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=1.92e-14 AS=2.24e-14 PD=5.6e-07 PS=6e-07 $X=106750 $Y=50125 $D=0
M1000 VDD 144 340 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 $X=107320 $Y=62980 $D=0
M1001 VDD 144 143 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 $X=107320 $Y=63840 $D=0
M1002 144 143 147 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=2.4e-14 AS=1.92e-14 PD=6.2e-07 PS=5.6e-07 $X=107320 $Y=64700 $D=0
M1003 147 141 144 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=2.4e-14 AS=2.4e-14 PD=6.2e-07 PS=6.2e-07 $X=107320 $Y=65100 $D=0
M1004 VDD 138 147 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=1.92e-14 AS=2.4e-14 PD=5.6e-07 PS=6.2e-07 $X=107320 $Y=65500 $D=0
M1005 VDD RESET 141 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 $X=107320 $Y=66360 $D=0
M1006 VDD 140 138 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 $X=107320 $Y=67220 $D=0
M1007 VDD CLK_MAIN 140 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 $X=107320 $Y=68080 $D=0
M1008 145 140 144 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 $X=107320 $Y=68940 $D=0
M1009 472 140 VDD VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=2.24e-14 AS=1.92e-14 PD=6e-07 PS=5.6e-07 $X=107320 $Y=69800 $D=0
M1010 142 145 472 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=1.92e-14 AS=2.24e-14 PD=5.6e-07 PS=6e-07 $X=107320 $Y=70180 $D=0
M1011 145 141 VDD VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=2.4e-14 AS=1.92e-14 PD=6.2e-07 PS=5.6e-07 $X=107320 $Y=71040 $D=0
M1012 VDD 142 145 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=1.92e-14 AS=2.4e-14 PD=5.6e-07 PS=6.2e-07 $X=107320 $Y=71440 $D=0
M1013 352 138 142 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 $X=107320 $Y=72300 $D=0
M1014 VDD 353 352 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 $X=107320 $Y=73160 $D=0
M1015 VDD B4 353 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 $X=107320 $Y=74020 $D=0
M1016 139 135 VDD VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=2.4e-14 AS=1.92e-14 PD=6.2e-07 PS=5.6e-07 $X=107610 $Y=50125 $D=0
M1017 VDD 351 148 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 $X=107790 $Y=58455 $D=0
M1018 355 121 VDD VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=1.84e-14 AS=1.84e-14 PD=5.5e-07 PS=5.5e-07 $X=107820 $Y=56315 $D=0
M1019 VDD 146 139 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=1.92e-14 AS=2.4e-14 PD=5.6e-07 PS=6.2e-07 $X=108010 $Y=50125 $D=0
M1020 SC4 121 148 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=2.24e-14 AS=1.84e-14 PD=6e-07 PS=5.5e-07 $X=108590 $Y=56315 $D=0
M1021 150 350 VDD VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 $X=108685 $Y=55295 $D=0
M1022 356 134 146 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 $X=108870 $Y=50125 $D=0
M1023 150 355 SC4 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=1.84e-14 AS=2.24e-14 PD=5.5e-07 PS=6e-07 $X=108970 $Y=56315 $D=0
M1024 VDD 357 356 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 $X=109730 $Y=50125 $D=0
M1025 VDD SC4 357 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 $X=110590 $Y=50125 $D=0
M1026 VDD 153 S5 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 $X=111970 $Y=50125 $D=0
M1027 VDD 153 154 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 $X=112830 $Y=50125 $D=0
M1028 VDD 359 365 VDD PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=2.07e-14 PD=6.4e-07 PS=5.9e-07 $X=113260 $Y=55725 $D=0
M1029 VDD 359 367 VDD PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=2.07e-14 PD=6.4e-07 PS=5.9e-07 $X=113260 $Y=58805 $D=0
M1030 VDD 360 359 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 $X=113515 $Y=61795 $D=0
M1031 VDD 158 360 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 $X=113525 $Y=62980 $D=0
M1032 VDD 158 157 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 $X=113525 $Y=63840 $D=0
M1033 158 157 161 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=2.4e-14 AS=1.92e-14 PD=6.2e-07 PS=5.6e-07 $X=113525 $Y=64700 $D=0
M1034 161 155 158 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=2.4e-14 AS=2.4e-14 PD=6.2e-07 PS=6.2e-07 $X=113525 $Y=65100 $D=0
M1035 VDD 151 161 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=1.92e-14 AS=2.4e-14 PD=5.6e-07 PS=6.2e-07 $X=113525 $Y=65500 $D=0
M1036 VDD RESET 155 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 $X=113525 $Y=66360 $D=0
M1037 VDD 152 151 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 $X=113525 $Y=67220 $D=0
M1038 VDD CLK_MAIN 152 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 $X=113525 $Y=68080 $D=0
M1039 159 152 158 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 $X=113525 $Y=68940 $D=0
M1040 473 152 VDD VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=2.24e-14 AS=1.92e-14 PD=6e-07 PS=5.6e-07 $X=113525 $Y=69800 $D=0
M1041 156 159 473 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=1.92e-14 AS=2.24e-14 PD=5.6e-07 PS=6e-07 $X=113525 $Y=70180 $D=0
M1042 159 155 VDD VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=2.4e-14 AS=1.92e-14 PD=6.2e-07 PS=5.6e-07 $X=113525 $Y=71040 $D=0
M1043 VDD 156 159 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=1.92e-14 AS=2.4e-14 PD=5.6e-07 PS=6.2e-07 $X=113525 $Y=71440 $D=0
M1044 361 151 156 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 $X=113525 $Y=72300 $D=0
M1045 VDD 362 361 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 $X=113525 $Y=73160 $D=0
M1046 VDD A5 362 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 $X=113525 $Y=74020 $D=0
M1047 365 363 VDD VDD PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=2.52e-14 PD=6.4e-07 PS=6.4e-07 $X=113640 $Y=55725 $D=0
M1048 367 363 VDD VDD PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=2.52e-14 PD=6.4e-07 PS=6.4e-07 $X=113640 $Y=58805 $D=0
M1049 153 154 160 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=2.4e-14 AS=1.92e-14 PD=6.2e-07 PS=5.6e-07 $X=113690 $Y=50125 $D=0
M1050 165 136 365 VDD PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=2.52e-14 PD=6.4e-07 PS=6.4e-07 $X=114020 $Y=55725 $D=0
M1051 166 137 367 VDD PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=2.52e-14 PD=6.4e-07 PS=6.4e-07 $X=114020 $Y=58805 $D=0
M1052 160 164 153 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=2.4e-14 AS=2.4e-14 PD=6.2e-07 PS=6.2e-07 $X=114090 $Y=50125 $D=0
M1053 474 359 165 VDD PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=2.52e-14 PD=6.4e-07 PS=6.4e-07 $X=114400 $Y=55725 $D=0
M1054 475 359 166 VDD PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=2.52e-14 PD=6.4e-07 PS=6.4e-07 $X=114400 $Y=58805 $D=0
M1055 VDD 163 160 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=1.92e-14 AS=2.4e-14 PD=5.6e-07 PS=6.2e-07 $X=114490 $Y=50125 $D=0
M1056 VDD 363 474 VDD PMOS_VTL L=5e-08 W=1.8e-07 AD=2.07e-14 AS=2.52e-14 PD=5.9e-07 PS=6.4e-07 $X=114780 $Y=55725 $D=0
M1057 VDD 363 475 VDD PMOS_VTL L=5e-08 W=1.8e-07 AD=2.07e-14 AS=2.52e-14 PD=5.9e-07 PS=6.4e-07 $X=114780 $Y=58805 $D=0
M1058 VDD RESET 164 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 $X=115350 $Y=50125 $D=0
M1059 370 359 VDD VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=2.24e-14 AS=1.84e-14 PD=6e-07 PS=5.5e-07 $X=115500 $Y=55725 $D=0
M1060 372 359 VDD VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=2.24e-14 AS=1.84e-14 PD=6e-07 PS=5.5e-07 $X=115500 $Y=58805 $D=0
M1061 VDD 363 370 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=2.24e-14 AS=2.24e-14 PD=6e-07 PS=6e-07 $X=115880 $Y=55725 $D=0
M1062 VDD 363 372 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=2.24e-14 AS=2.24e-14 PD=6e-07 PS=6e-07 $X=115880 $Y=58805 $D=0
M1063 VDD 162 163 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 $X=116210 $Y=50125 $D=0
M1064 370 136 VDD VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=1.84e-14 AS=2.24e-14 PD=5.5e-07 PS=6e-07 $X=116260 $Y=55725 $D=0
M1065 372 137 VDD VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=1.84e-14 AS=2.24e-14 PD=5.5e-07 PS=6e-07 $X=116260 $Y=58805 $D=0
M1066 179 165 370 VDD PMOS_VTL L=5e-08 W=1.4e-07 AD=1.68e-14 AS=1.75e-14 PD=5.2e-07 PS=5.3e-07 $X=117000 $Y=55725 $D=0
M1067 177 166 372 VDD PMOS_VTL L=5e-08 W=1.4e-07 AD=1.68e-14 AS=1.75e-14 PD=5.2e-07 PS=5.3e-07 $X=117000 $Y=58805 $D=0
M1068 VDD CLK_MAIN 162 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 $X=117070 $Y=50125 $D=0
M1069 476 136 179 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=2.24e-14 AS=1.84e-14 PD=6e-07 PS=5.5e-07 $X=117730 $Y=55725 $D=0
M1070 477 137 177 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=2.24e-14 AS=1.84e-14 PD=6e-07 PS=5.5e-07 $X=117730 $Y=58805 $D=0
M1071 169 162 153 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 $X=117930 $Y=50125 $D=0
M1072 478 359 476 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=2.24e-14 AS=2.24e-14 PD=6e-07 PS=6e-07 $X=118110 $Y=55725 $D=0
M1073 479 359 477 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=2.24e-14 AS=2.24e-14 PD=6e-07 PS=6e-07 $X=118110 $Y=58805 $D=0
M1074 VDD 363 478 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=1.84e-14 AS=2.24e-14 PD=5.5e-07 PS=6e-07 $X=118490 $Y=55725 $D=0
M1075 VDD 363 479 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=1.84e-14 AS=2.24e-14 PD=5.5e-07 PS=6e-07 $X=118490 $Y=58805 $D=0
M1076 480 162 VDD VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=2.24e-14 AS=1.92e-14 PD=6e-07 PS=5.6e-07 $X=118790 $Y=50125 $D=0
M1077 VDD 373 363 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 $X=119035 $Y=61795 $D=0
M1078 VDD 173 373 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 $X=119045 $Y=62980 $D=0
M1079 VDD 173 172 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 $X=119045 $Y=63840 $D=0
M1080 173 172 175 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=2.4e-14 AS=1.92e-14 PD=6.2e-07 PS=5.6e-07 $X=119045 $Y=64700 $D=0
M1081 175 170 173 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=2.4e-14 AS=2.4e-14 PD=6.2e-07 PS=6.2e-07 $X=119045 $Y=65100 $D=0
M1082 VDD 167 175 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=1.92e-14 AS=2.4e-14 PD=5.6e-07 PS=6.2e-07 $X=119045 $Y=65500 $D=0
M1083 VDD RESET 170 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 $X=119045 $Y=66360 $D=0
M1084 VDD 168 167 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 $X=119045 $Y=67220 $D=0
M1085 VDD CLK_MAIN 168 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 $X=119045 $Y=68080 $D=0
M1086 174 168 173 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 $X=119045 $Y=68940 $D=0
M1087 481 168 VDD VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=2.24e-14 AS=1.92e-14 PD=6e-07 PS=5.6e-07 $X=119045 $Y=69800 $D=0
M1088 171 174 481 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=1.92e-14 AS=2.24e-14 PD=5.6e-07 PS=6e-07 $X=119045 $Y=70180 $D=0
M1089 174 170 VDD VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=2.4e-14 AS=1.92e-14 PD=6.2e-07 PS=5.6e-07 $X=119045 $Y=71040 $D=0
M1090 VDD 171 174 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=1.92e-14 AS=2.4e-14 PD=5.6e-07 PS=6.2e-07 $X=119045 $Y=71440 $D=0
M1091 374 167 171 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 $X=119045 $Y=72300 $D=0
M1092 VDD 375 374 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 $X=119045 $Y=73160 $D=0
M1093 VDD B5 375 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 $X=119045 $Y=74020 $D=0
M1094 176 169 480 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=1.92e-14 AS=2.24e-14 PD=5.6e-07 PS=6e-07 $X=119170 $Y=50125 $D=0
M1095 377 121 VDD VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=1.84e-14 AS=1.84e-14 PD=5.5e-07 PS=5.5e-07 $X=119620 $Y=56265 $D=0
M1096 169 164 VDD VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=2.4e-14 AS=1.92e-14 PD=6.2e-07 PS=5.6e-07 $X=120030 $Y=50125 $D=0
M1097 SC5 121 177 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=2.24e-14 AS=1.84e-14 PD=6e-07 PS=5.5e-07 $X=120390 $Y=56265 $D=0
M1098 VDD 176 169 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=1.92e-14 AS=2.4e-14 PD=5.6e-07 PS=6.2e-07 $X=120430 $Y=50125 $D=0
M1099 179 377 SC5 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=1.84e-14 AS=2.24e-14 PD=5.5e-07 PS=6e-07 $X=120770 $Y=56265 $D=0
M1100 378 163 176 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 $X=121290 $Y=50125 $D=0
M1101 VDD 379 378 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 $X=122150 $Y=50125 $D=0
M1102 VDD SC5 379 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 $X=123010 $Y=50125 $D=0
M1103 VDD 182 S6 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 $X=124525 $Y=50125 $D=0
M1104 VDD 381 386 VDD PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=2.07e-14 PD=6.4e-07 PS=5.9e-07 $X=125060 $Y=55775 $D=0
M1105 VDD 381 388 VDD PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=2.07e-14 PD=6.4e-07 PS=5.9e-07 $X=125060 $Y=58855 $D=0
M1106 VDD 182 185 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 $X=125385 $Y=50125 $D=0
M1107 VDD 187 381 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 $X=125420 $Y=62980 $D=0
M1108 VDD 187 186 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 $X=125420 $Y=63840 $D=0
M1109 187 186 189 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=2.4e-14 AS=1.92e-14 PD=6.2e-07 PS=5.6e-07 $X=125420 $Y=64700 $D=0
M1110 189 183 187 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=2.4e-14 AS=2.4e-14 PD=6.2e-07 PS=6.2e-07 $X=125420 $Y=65100 $D=0
M1111 VDD 180 189 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=1.92e-14 AS=2.4e-14 PD=5.6e-07 PS=6.2e-07 $X=125420 $Y=65500 $D=0
M1112 VDD RESET 183 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 $X=125420 $Y=66360 $D=0
M1113 VDD 181 180 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 $X=125420 $Y=67220 $D=0
M1114 VDD CLK_MAIN 181 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 $X=125420 $Y=68080 $D=0
M1115 188 181 187 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 $X=125420 $Y=68940 $D=0
M1116 482 181 VDD VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=2.24e-14 AS=1.92e-14 PD=6e-07 PS=5.6e-07 $X=125420 $Y=69800 $D=0
M1117 184 188 482 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=1.92e-14 AS=2.24e-14 PD=5.6e-07 PS=6e-07 $X=125420 $Y=70180 $D=0
M1118 188 183 VDD VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=2.4e-14 AS=1.92e-14 PD=6.2e-07 PS=5.6e-07 $X=125420 $Y=71040 $D=0
M1119 VDD 184 188 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=1.92e-14 AS=2.4e-14 PD=5.6e-07 PS=6.2e-07 $X=125420 $Y=71440 $D=0
M1120 382 180 184 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 $X=125420 $Y=72300 $D=0
M1121 VDD 383 382 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 $X=125420 $Y=73160 $D=0
M1122 VDD A6 383 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 $X=125420 $Y=74020 $D=0
M1123 386 384 VDD VDD PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=2.52e-14 PD=6.4e-07 PS=6.4e-07 $X=125440 $Y=55775 $D=0
M1124 388 384 VDD VDD PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=2.52e-14 PD=6.4e-07 PS=6.4e-07 $X=125440 $Y=58855 $D=0
M1125 194 165 386 VDD PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=2.52e-14 PD=6.4e-07 PS=6.4e-07 $X=125820 $Y=55775 $D=0
M1126 195 166 388 VDD PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=2.52e-14 PD=6.4e-07 PS=6.4e-07 $X=125820 $Y=58855 $D=0
M1127 483 381 194 VDD PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=2.52e-14 PD=6.4e-07 PS=6.4e-07 $X=126200 $Y=55775 $D=0
M1128 484 381 195 VDD PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=2.52e-14 PD=6.4e-07 PS=6.4e-07 $X=126200 $Y=58855 $D=0
M1129 182 185 190 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=2.4e-14 AS=1.92e-14 PD=6.2e-07 PS=5.6e-07 $X=126245 $Y=50125 $D=0
M1130 VDD 384 483 VDD PMOS_VTL L=5e-08 W=1.8e-07 AD=2.07e-14 AS=2.52e-14 PD=5.9e-07 PS=6.4e-07 $X=126580 $Y=55775 $D=0
M1131 VDD 384 484 VDD PMOS_VTL L=5e-08 W=1.8e-07 AD=2.07e-14 AS=2.52e-14 PD=5.9e-07 PS=6.4e-07 $X=126580 $Y=58855 $D=0
M1132 190 193 182 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=2.4e-14 AS=2.4e-14 PD=6.2e-07 PS=6.2e-07 $X=126645 $Y=50125 $D=0
M1133 VDD 192 190 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=1.92e-14 AS=2.4e-14 PD=5.6e-07 PS=6.2e-07 $X=127045 $Y=50125 $D=0
M1134 391 381 VDD VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=2.24e-14 AS=1.84e-14 PD=6e-07 PS=5.5e-07 $X=127300 $Y=55775 $D=0
M1135 393 381 VDD VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=2.24e-14 AS=1.84e-14 PD=6e-07 PS=5.5e-07 $X=127300 $Y=58855 $D=0
M1136 VDD 384 391 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=2.24e-14 AS=2.24e-14 PD=6e-07 PS=6e-07 $X=127680 $Y=55775 $D=0
M1137 VDD 384 393 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=2.24e-14 AS=2.24e-14 PD=6e-07 PS=6e-07 $X=127680 $Y=58855 $D=0
M1138 VDD RESET 193 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 $X=127905 $Y=50125 $D=0
M1139 391 165 VDD VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=1.84e-14 AS=2.24e-14 PD=5.5e-07 PS=6e-07 $X=128060 $Y=55775 $D=0
M1140 393 166 VDD VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=1.84e-14 AS=2.24e-14 PD=5.5e-07 PS=6e-07 $X=128060 $Y=58855 $D=0
M1141 VDD 191 192 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 $X=128765 $Y=50125 $D=0
M1142 394 194 391 VDD PMOS_VTL L=5e-08 W=1.4e-07 AD=1.68e-14 AS=1.75e-14 PD=5.2e-07 PS=5.3e-07 $X=128800 $Y=55775 $D=0
M1143 395 195 393 VDD PMOS_VTL L=5e-08 W=1.4e-07 AD=1.68e-14 AS=1.75e-14 PD=5.2e-07 PS=5.3e-07 $X=128800 $Y=58855 $D=0
M1144 485 165 394 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=2.24e-14 AS=1.84e-14 PD=6e-07 PS=5.5e-07 $X=129530 $Y=55775 $D=0
M1145 486 166 395 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=2.24e-14 AS=1.84e-14 PD=6e-07 PS=5.5e-07 $X=129530 $Y=58855 $D=0
M1146 VDD CLK_MAIN 191 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 $X=129625 $Y=50125 $D=0
M1147 487 381 485 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=2.24e-14 AS=2.24e-14 PD=6e-07 PS=6e-07 $X=129910 $Y=55775 $D=0
M1148 488 381 486 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=2.24e-14 AS=2.24e-14 PD=6e-07 PS=6e-07 $X=129910 $Y=58855 $D=0
M1149 VDD 384 487 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=1.84e-14 AS=2.24e-14 PD=5.5e-07 PS=6e-07 $X=130290 $Y=55775 $D=0
M1150 VDD 384 488 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=1.84e-14 AS=2.24e-14 PD=5.5e-07 PS=6e-07 $X=130290 $Y=58855 $D=0
M1151 203 191 182 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 $X=130485 $Y=50125 $D=0
M1152 VDD 201 384 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 $X=130920 $Y=62980 $D=0
M1153 VDD 201 200 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 $X=130920 $Y=63840 $D=0
M1154 201 200 204 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=2.4e-14 AS=1.92e-14 PD=6.2e-07 PS=5.6e-07 $X=130920 $Y=64700 $D=0
M1155 204 198 201 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=2.4e-14 AS=2.4e-14 PD=6.2e-07 PS=6.2e-07 $X=130920 $Y=65100 $D=0
M1156 VDD 196 204 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=1.92e-14 AS=2.4e-14 PD=5.6e-07 PS=6.2e-07 $X=130920 $Y=65500 $D=0
M1157 VDD RESET 198 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 $X=130920 $Y=66360 $D=0
M1158 VDD 197 196 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 $X=130920 $Y=67220 $D=0
M1159 VDD CLK_MAIN 197 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 $X=130920 $Y=68080 $D=0
M1160 202 197 201 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 $X=130920 $Y=68940 $D=0
M1161 489 197 VDD VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=2.24e-14 AS=1.92e-14 PD=6e-07 PS=5.6e-07 $X=130920 $Y=69800 $D=0
M1162 199 202 489 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=1.92e-14 AS=2.24e-14 PD=5.6e-07 PS=6e-07 $X=130920 $Y=70180 $D=0
M1163 202 198 VDD VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=2.4e-14 AS=1.92e-14 PD=6.2e-07 PS=5.6e-07 $X=130920 $Y=71040 $D=0
M1164 VDD 199 202 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=1.92e-14 AS=2.4e-14 PD=5.6e-07 PS=6.2e-07 $X=130920 $Y=71440 $D=0
M1165 396 196 199 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 $X=130920 $Y=72300 $D=0
M1166 VDD 397 396 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 $X=130920 $Y=73160 $D=0
M1167 VDD B6 397 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 $X=130920 $Y=74020 $D=0
M1168 490 191 VDD VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=2.24e-14 AS=1.92e-14 PD=6e-07 PS=5.6e-07 $X=131345 $Y=50125 $D=0
M1169 VDD 395 206 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 $X=131390 $Y=58455 $D=0
M1170 399 121 VDD VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=1.84e-14 AS=1.84e-14 PD=5.5e-07 PS=5.5e-07 $X=131420 $Y=56315 $D=0
M1171 205 203 490 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=1.92e-14 AS=2.24e-14 PD=5.6e-07 PS=6e-07 $X=131725 $Y=50125 $D=0
M1172 SC6 121 206 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=2.24e-14 AS=1.84e-14 PD=6e-07 PS=5.5e-07 $X=132190 $Y=56315 $D=0
M1173 208 394 VDD VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 $X=132285 $Y=55135 $D=0
M1174 208 399 SC6 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=1.84e-14 AS=2.24e-14 PD=5.5e-07 PS=6e-07 $X=132570 $Y=56315 $D=0
M1175 203 193 VDD VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=2.4e-14 AS=1.92e-14 PD=6.2e-07 PS=5.6e-07 $X=132585 $Y=50125 $D=0
M1176 VDD 205 203 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=1.92e-14 AS=2.4e-14 PD=5.6e-07 PS=6.2e-07 $X=132985 $Y=50125 $D=0
M1177 400 192 205 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 $X=133845 $Y=50125 $D=0
M1178 VDD 401 400 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 $X=134705 $Y=50125 $D=0
M1179 VDD SC6 401 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 $X=135565 $Y=50125 $D=0
M1180 VDD 403 409 VDD PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=2.07e-14 PD=6.4e-07 PS=5.9e-07 $X=136860 $Y=55775 $D=0
M1181 VDD 403 411 VDD PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=2.07e-14 PD=6.4e-07 PS=5.9e-07 $X=136860 $Y=58855 $D=0
M1182 VDD 216 S7 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 $X=136905 $Y=50125 $D=0
M1183 VDD 404 403 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 $X=137115 $Y=61795 $D=0
M1184 VDD 214 404 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 $X=137125 $Y=62980 $D=0
M1185 VDD 214 213 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 $X=137125 $Y=63840 $D=0
M1186 214 213 217 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=2.4e-14 AS=1.92e-14 PD=6.2e-07 PS=5.6e-07 $X=137125 $Y=64700 $D=0
M1187 217 211 214 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=2.4e-14 AS=2.4e-14 PD=6.2e-07 PS=6.2e-07 $X=137125 $Y=65100 $D=0
M1188 VDD 209 217 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=1.92e-14 AS=2.4e-14 PD=5.6e-07 PS=6.2e-07 $X=137125 $Y=65500 $D=0
M1189 VDD RESET 211 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 $X=137125 $Y=66360 $D=0
M1190 VDD 210 209 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 $X=137125 $Y=67220 $D=0
M1191 VDD CLK_MAIN 210 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 $X=137125 $Y=68080 $D=0
M1192 215 210 214 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 $X=137125 $Y=68940 $D=0
M1193 491 210 VDD VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=2.24e-14 AS=1.92e-14 PD=6e-07 PS=5.6e-07 $X=137125 $Y=69800 $D=0
M1194 212 215 491 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=1.92e-14 AS=2.24e-14 PD=5.6e-07 PS=6e-07 $X=137125 $Y=70180 $D=0
M1195 215 211 VDD VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=2.4e-14 AS=1.92e-14 PD=6.2e-07 PS=5.6e-07 $X=137125 $Y=71040 $D=0
M1196 VDD 212 215 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=1.92e-14 AS=2.4e-14 PD=5.6e-07 PS=6.2e-07 $X=137125 $Y=71440 $D=0
M1197 405 209 212 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 $X=137125 $Y=72300 $D=0
M1198 VDD 406 405 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 $X=137125 $Y=73160 $D=0
M1199 VDD A7 406 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 $X=137125 $Y=74020 $D=0
M1200 409 407 VDD VDD PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=2.52e-14 PD=6.4e-07 PS=6.4e-07 $X=137240 $Y=55775 $D=0
M1201 411 407 VDD VDD PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=2.52e-14 PD=6.4e-07 PS=6.4e-07 $X=137240 $Y=58855 $D=0
M1202 223 194 409 VDD PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=2.52e-14 PD=6.4e-07 PS=6.4e-07 $X=137620 $Y=55775 $D=0
M1203 224 195 411 VDD PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=2.52e-14 PD=6.4e-07 PS=6.4e-07 $X=137620 $Y=58855 $D=0
M1204 VDD 216 218 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 $X=137765 $Y=50125 $D=0
M1205 492 403 223 VDD PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=2.52e-14 PD=6.4e-07 PS=6.4e-07 $X=138000 $Y=55775 $D=0
M1206 493 403 224 VDD PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=2.52e-14 PD=6.4e-07 PS=6.4e-07 $X=138000 $Y=58855 $D=0
M1207 VDD 407 492 VDD PMOS_VTL L=5e-08 W=1.8e-07 AD=2.07e-14 AS=2.52e-14 PD=5.9e-07 PS=6.4e-07 $X=138380 $Y=55775 $D=0
M1208 VDD 407 493 VDD PMOS_VTL L=5e-08 W=1.8e-07 AD=2.07e-14 AS=2.52e-14 PD=5.9e-07 PS=6.4e-07 $X=138380 $Y=58855 $D=0
M1209 216 218 219 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=2.4e-14 AS=1.92e-14 PD=6.2e-07 PS=5.6e-07 $X=138625 $Y=50125 $D=0
M1210 219 222 216 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=2.4e-14 AS=2.4e-14 PD=6.2e-07 PS=6.2e-07 $X=139025 $Y=50125 $D=0
M1211 414 403 VDD VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=2.24e-14 AS=1.84e-14 PD=6e-07 PS=5.5e-07 $X=139100 $Y=55775 $D=0
M1212 416 403 VDD VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=2.24e-14 AS=1.84e-14 PD=6e-07 PS=5.5e-07 $X=139100 $Y=58855 $D=0
M1213 VDD 221 219 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=1.92e-14 AS=2.4e-14 PD=5.6e-07 PS=6.2e-07 $X=139425 $Y=50125 $D=0
M1214 VDD 407 414 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=2.24e-14 AS=2.24e-14 PD=6e-07 PS=6e-07 $X=139480 $Y=55775 $D=0
M1215 VDD 407 416 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=2.24e-14 AS=2.24e-14 PD=6e-07 PS=6e-07 $X=139480 $Y=58855 $D=0
M1216 414 194 VDD VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=1.84e-14 AS=2.24e-14 PD=5.5e-07 PS=6e-07 $X=139860 $Y=55775 $D=0
M1217 416 195 VDD VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=1.84e-14 AS=2.24e-14 PD=5.5e-07 PS=6e-07 $X=139860 $Y=58855 $D=0
M1218 VDD RESET 222 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 $X=140285 $Y=50125 $D=0
M1219 237 223 414 VDD PMOS_VTL L=5e-08 W=1.4e-07 AD=1.68e-14 AS=1.75e-14 PD=5.2e-07 PS=5.3e-07 $X=140600 $Y=55775 $D=0
M1220 234 224 416 VDD PMOS_VTL L=5e-08 W=1.4e-07 AD=1.68e-14 AS=1.75e-14 PD=5.2e-07 PS=5.3e-07 $X=140600 $Y=58855 $D=0
M1221 VDD 220 221 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 $X=141145 $Y=50125 $D=0
M1222 494 194 237 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=2.24e-14 AS=1.84e-14 PD=6e-07 PS=5.5e-07 $X=141330 $Y=55775 $D=0
M1223 495 195 234 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=2.24e-14 AS=1.84e-14 PD=6e-07 PS=5.5e-07 $X=141330 $Y=58855 $D=0
M1224 496 403 494 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=2.24e-14 AS=2.24e-14 PD=6e-07 PS=6e-07 $X=141710 $Y=55775 $D=0
M1225 497 403 495 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=2.24e-14 AS=2.24e-14 PD=6e-07 PS=6e-07 $X=141710 $Y=58855 $D=0
M1226 VDD CLK_MAIN 220 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 $X=142005 $Y=50125 $D=0
M1227 VDD 407 496 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=1.84e-14 AS=2.24e-14 PD=5.5e-07 PS=6e-07 $X=142090 $Y=55775 $D=0
M1228 VDD 407 497 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=1.84e-14 AS=2.24e-14 PD=5.5e-07 PS=6e-07 $X=142090 $Y=58855 $D=0
M1229 VDD 417 407 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 $X=142635 $Y=61795 $D=0
M1230 VDD 230 417 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 $X=142645 $Y=62980 $D=0
M1231 VDD 230 229 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 $X=142645 $Y=63840 $D=0
M1232 230 229 232 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=2.4e-14 AS=1.92e-14 PD=6.2e-07 PS=5.6e-07 $X=142645 $Y=64700 $D=0
M1233 232 227 230 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=2.4e-14 AS=2.4e-14 PD=6.2e-07 PS=6.2e-07 $X=142645 $Y=65100 $D=0
M1234 VDD 225 232 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=1.92e-14 AS=2.4e-14 PD=5.6e-07 PS=6.2e-07 $X=142645 $Y=65500 $D=0
M1235 VDD RESET 227 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 $X=142645 $Y=66360 $D=0
M1236 VDD 226 225 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 $X=142645 $Y=67220 $D=0
M1237 VDD CLK_MAIN 226 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 $X=142645 $Y=68080 $D=0
M1238 231 226 230 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 $X=142645 $Y=68940 $D=0
M1239 498 226 VDD VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=2.24e-14 AS=1.92e-14 PD=6e-07 PS=5.6e-07 $X=142645 $Y=69800 $D=0
M1240 228 231 498 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=1.92e-14 AS=2.24e-14 PD=5.6e-07 PS=6e-07 $X=142645 $Y=70180 $D=0
M1241 231 227 VDD VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=2.4e-14 AS=1.92e-14 PD=6.2e-07 PS=5.6e-07 $X=142645 $Y=71040 $D=0
M1242 VDD 228 231 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=1.92e-14 AS=2.4e-14 PD=5.6e-07 PS=6.2e-07 $X=142645 $Y=71440 $D=0
M1243 418 225 228 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 $X=142645 $Y=72300 $D=0
M1244 VDD 419 418 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 $X=142645 $Y=73160 $D=0
M1245 VDD B7 419 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 $X=142645 $Y=74020 $D=0
M1246 233 220 216 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 $X=142865 $Y=50125 $D=0
M1247 421 121 VDD VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=1.84e-14 AS=1.84e-14 PD=5.5e-07 PS=5.5e-07 $X=143220 $Y=56315 $D=0
M1248 499 220 VDD VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=2.24e-14 AS=1.92e-14 PD=6e-07 PS=5.6e-07 $X=143725 $Y=50125 $D=0
M1249 SC7 121 234 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=2.24e-14 AS=1.84e-14 PD=6e-07 PS=5.5e-07 $X=143990 $Y=56315 $D=0
M1250 236 233 499 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=1.92e-14 AS=2.24e-14 PD=5.6e-07 PS=6e-07 $X=144105 $Y=50125 $D=0
M1251 237 421 SC7 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=1.84e-14 AS=2.24e-14 PD=5.5e-07 PS=6e-07 $X=144370 $Y=56315 $D=0
M1252 233 222 VDD VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=2.4e-14 AS=1.92e-14 PD=6.2e-07 PS=5.6e-07 $X=144965 $Y=50125 $D=0
M1253 VDD 236 233 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=1.92e-14 AS=2.4e-14 PD=5.6e-07 PS=6.2e-07 $X=145365 $Y=50125 $D=0
M1254 423 221 236 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 $X=146225 $Y=50125 $D=0
M1255 422 121 VDD VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=1.84e-14 AS=1.84e-14 PD=5.5e-07 PS=5.5e-07 $X=146325 $Y=56290 $D=0
M1256 VDD 424 423 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 $X=147085 $Y=50125 $D=0
M1257 C7_OUT 121 224 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=2.24e-14 AS=1.84e-14 PD=6e-07 PS=5.5e-07 $X=147095 $Y=56290 $D=0
M1258 223 422 C7_OUT VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=1.84e-14 AS=2.24e-14 PD=5.5e-07 PS=6e-07 $X=147475 $Y=56290 $D=0
M1259 VDD SC7 424 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 $X=147945 $Y=50125 $D=0
M1260 426 C7_OUT VDD VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 $X=149095 $Y=57685 $D=0
M1261 427 426 VDD VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 $X=149095 $Y=58545 $D=0
M1262 245 239 427 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 $X=149095 $Y=59405 $D=0
M1263 246 245 VDD VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=2.4e-14 AS=1.92e-14 PD=6.2e-07 PS=5.6e-07 $X=149095 $Y=60265 $D=0
M1264 VDD 242 246 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=1.92e-14 AS=2.4e-14 PD=5.6e-07 PS=6.2e-07 $X=149095 $Y=60665 $D=0
M1265 500 246 245 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=2.24e-14 AS=1.92e-14 PD=6e-07 PS=5.6e-07 $X=149095 $Y=61525 $D=0
M1266 VDD 243 500 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=1.92e-14 AS=2.24e-14 PD=5.6e-07 PS=6e-07 $X=149095 $Y=61905 $D=0
M1267 241 243 246 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 $X=149095 $Y=62765 $D=0
M1268 243 CLK_MAIN VDD VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 $X=149095 $Y=63625 $D=0
M1269 239 243 VDD VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 $X=149095 $Y=64485 $D=0
M1270 242 RESET VDD VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 $X=149095 $Y=65345 $D=0
M1271 244 239 VDD VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=2.4e-14 AS=1.92e-14 PD=6.2e-07 PS=5.6e-07 $X=149095 $Y=66205 $D=0
M1272 241 242 244 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=2.4e-14 AS=2.4e-14 PD=6.2e-07 PS=6.2e-07 $X=149095 $Y=66605 $D=0
M1273 244 240 241 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=1.92e-14 AS=2.4e-14 PD=5.6e-07 PS=6.2e-07 $X=149095 $Y=67005 $D=0
M1274 240 241 VDD VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 $X=149095 $Y=67865 $D=0
M1275 Cout 241 VDD VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 $X=149095 $Y=68725 $D=0
.ENDS
***************************************
