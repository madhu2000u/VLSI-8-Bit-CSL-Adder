* SPICE NETLIST
***************************************

.SUBCKT 1_bit_mirror_full_adder A B Cin ~Cout ~S GND VDD
** N=17 EP=7 IP=0 FDC=24
M0 GND A 3 GND NMOS_VTL L=5e-08 W=2.7e-07 AD=3.78e-14 AS=3.105e-14 PD=8.2e-07 PS=7.7e-07 $X=81449430 $Y=33694290 $D=1
M1 3 B GND GND NMOS_VTL L=5e-08 W=2.7e-07 AD=3.78e-14 AS=3.78e-14 PD=8.2e-07 PS=8.2e-07 $X=81449810 $Y=33694290 $D=1
M2 ~Cout Cin 3 GND NMOS_VTL L=5e-08 W=2.7e-07 AD=3.78e-14 AS=3.78e-14 PD=8.2e-07 PS=8.2e-07 $X=81450190 $Y=33694290 $D=1
M3 15 A ~Cout GND NMOS_VTL L=5e-08 W=2.7e-07 AD=3.78e-14 AS=3.78e-14 PD=8.2e-07 PS=8.2e-07 $X=81450570 $Y=33694290 $D=1
M4 GND B 15 GND NMOS_VTL L=5e-08 W=2.7e-07 AD=3.105e-14 AS=3.78e-14 PD=7.7e-07 PS=8.2e-07 $X=81450950 $Y=33694290 $D=1
M5 7 A GND GND NMOS_VTL L=5e-08 W=2.7e-07 AD=3.78e-14 AS=3.105e-14 PD=8.2e-07 PS=7.7e-07 $X=81451670 $Y=33694290 $D=1
M6 GND B 7 GND NMOS_VTL L=5e-08 W=2.7e-07 AD=3.78e-14 AS=3.78e-14 PD=8.2e-07 PS=8.2e-07 $X=81452050 $Y=33694290 $D=1
M7 7 Cin GND GND NMOS_VTL L=5e-08 W=2.7e-07 AD=3.105e-14 AS=3.78e-14 PD=7.7e-07 PS=8.2e-07 $X=81452430 $Y=33694290 $D=1
M8 ~S ~Cout 7 GND NMOS_VTL L=5e-08 W=2.7e-07 AD=3.24e-14 AS=3.375e-14 PD=7.8e-07 PS=7.9e-07 $X=81453170 $Y=33694290 $D=1
M9 16 Cin ~S GND NMOS_VTL L=5e-08 W=2.7e-07 AD=3.78e-14 AS=3.105e-14 PD=8.2e-07 PS=7.7e-07 $X=81453900 $Y=33694290 $D=1
M10 17 A 16 GND NMOS_VTL L=5e-08 W=2.7e-07 AD=3.78e-14 AS=3.78e-14 PD=8.2e-07 PS=8.2e-07 $X=81454280 $Y=33694290 $D=1
M11 GND B 17 GND NMOS_VTL L=5e-08 W=2.7e-07 AD=3.105e-14 AS=3.78e-14 PD=7.7e-07 PS=8.2e-07 $X=81454660 $Y=33694290 $D=1
M12 VDD A 4 VDD PMOS_VTL L=5e-08 W=4e-07 AD=5.6e-14 AS=4.6e-14 PD=1.08e-06 PS=1.03e-06 $X=81449430 $Y=33695810 $D=0
M13 4 B VDD VDD PMOS_VTL L=5e-08 W=4e-07 AD=5.6e-14 AS=5.6e-14 PD=1.08e-06 PS=1.08e-06 $X=81449810 $Y=33695810 $D=0
M14 ~Cout Cin 4 VDD PMOS_VTL L=5e-08 W=4e-07 AD=5.6e-14 AS=5.6e-14 PD=1.08e-06 PS=1.08e-06 $X=81450190 $Y=33695810 $D=0
M15 12 A ~Cout VDD PMOS_VTL L=5e-08 W=4e-07 AD=5.6e-14 AS=5.6e-14 PD=1.08e-06 PS=1.08e-06 $X=81450570 $Y=33695810 $D=0
M16 VDD B 12 VDD PMOS_VTL L=5e-08 W=4e-07 AD=4.6e-14 AS=5.6e-14 PD=1.03e-06 PS=1.08e-06 $X=81450950 $Y=33695810 $D=0
M17 8 A VDD VDD PMOS_VTL L=5e-08 W=4e-07 AD=5.6e-14 AS=4.6e-14 PD=1.08e-06 PS=1.03e-06 $X=81451670 $Y=33695810 $D=0
M18 VDD B 8 VDD PMOS_VTL L=5e-08 W=4e-07 AD=5.6e-14 AS=5.6e-14 PD=1.08e-06 PS=1.08e-06 $X=81452050 $Y=33695810 $D=0
M19 8 Cin VDD VDD PMOS_VTL L=5e-08 W=4e-07 AD=4.6e-14 AS=5.6e-14 PD=1.03e-06 PS=1.08e-06 $X=81452430 $Y=33695810 $D=0
M20 ~S ~Cout 8 VDD PMOS_VTL L=5e-08 W=4e-07 AD=4.8e-14 AS=5e-14 PD=1.04e-06 PS=1.05e-06 $X=81453170 $Y=33695810 $D=0
M21 13 Cin ~S VDD PMOS_VTL L=5e-08 W=4e-07 AD=5.6e-14 AS=4.6e-14 PD=1.08e-06 PS=1.03e-06 $X=81453900 $Y=33695810 $D=0
M22 14 A 13 VDD PMOS_VTL L=5e-08 W=4e-07 AD=5.6e-14 AS=5.6e-14 PD=1.08e-06 PS=1.08e-06 $X=81454280 $Y=33695810 $D=0
M23 VDD B 14 VDD PMOS_VTL L=5e-08 W=4e-07 AD=4.6e-14 AS=5.6e-14 PD=1.03e-06 PS=1.08e-06 $X=81454660 $Y=33695810 $D=0
.ENDS
***************************************
