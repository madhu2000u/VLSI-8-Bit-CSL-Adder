/home/home5/msudhanan/ese555workingdir/sim_8_Bit_CSL_Adder_svrun1/ihnl/cds1/netlist