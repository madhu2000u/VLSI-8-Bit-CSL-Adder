* SPICE NETLIST
***************************************

.SUBCKT D_flip_flop D CLK_MAIN RESET GND VDD Q
** N=21 EP=6 IP=0 FDC=32
M0 10 D GND GND NMOS_VTL L=5e-08 W=1e-07 AD=1.2e-14 AS=1.2e-14 PD=4.4e-07 PS=4.4e-07 $X=4040 $Y=980 $D=1
M1 11 10 GND GND NMOS_VTL L=5e-08 W=1e-07 AD=1.2e-14 AS=1.2e-14 PD=4.4e-07 PS=4.4e-07 $X=4900 $Y=980 $D=1
M2 3 1 11 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.2e-14 AS=1.2e-14 PD=4.4e-07 PS=4.4e-07 $X=5760 $Y=980 $D=1
M3 18 3 GND GND NMOS_VTL L=5e-08 W=1e-07 AD=1.5e-14 AS=1.2e-14 PD=5e-07 PS=4.4e-07 $X=6620 $Y=980 $D=1
M4 5 4 18 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.2e-14 AS=1.5e-14 PD=4.4e-07 PS=5e-07 $X=7020 $Y=980 $D=1
M5 19 5 3 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.4e-14 AS=1.2e-14 PD=4.8e-07 PS=4.4e-07 $X=7880 $Y=980 $D=1
M6 GND 2 19 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.2e-14 AS=1.4e-14 PD=4.4e-07 PS=4.8e-07 $X=8260 $Y=980 $D=1
M7 6 2 5 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.2e-14 AS=1.2e-14 PD=4.4e-07 PS=4.4e-07 $X=9120 $Y=980 $D=1
M8 1 CLK_MAIN GND GND NMOS_VTL L=5e-08 W=1e-07 AD=1.2e-14 AS=1.2e-14 PD=4.4e-07 PS=4.4e-07 $X=9980 $Y=980 $D=1
M9 2 1 GND GND NMOS_VTL L=5e-08 W=1e-07 AD=1.2e-14 AS=1.2e-14 PD=4.4e-07 PS=4.4e-07 $X=10840 $Y=980 $D=1
M10 4 RESET GND GND NMOS_VTL L=5e-08 W=1e-07 AD=1.2e-14 AS=1.2e-14 PD=4.4e-07 PS=4.4e-07 $X=11700 $Y=980 $D=1
M11 20 1 GND GND NMOS_VTL L=5e-08 W=1e-07 AD=1.4e-14 AS=1.2e-14 PD=4.8e-07 PS=4.4e-07 $X=12580 $Y=980 $D=1
M12 21 4 20 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.5e-14 AS=1.4e-14 PD=5e-07 PS=4.8e-07 $X=12960 $Y=980 $D=1
M13 6 8 21 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.2e-14 AS=1.5e-14 PD=4.4e-07 PS=5e-07 $X=13360 $Y=980 $D=1
M14 8 6 GND GND NMOS_VTL L=5e-08 W=1e-07 AD=1.2e-14 AS=1.2e-14 PD=4.4e-07 PS=4.4e-07 $X=14220 $Y=980 $D=1
M15 Q 6 GND GND NMOS_VTL L=5e-08 W=1e-07 AD=1.2e-14 AS=1.2e-14 PD=4.4e-07 PS=4.4e-07 $X=15080 $Y=980 $D=1
M16 10 D VDD VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 $X=4040 $Y=1880 $D=0
M17 11 10 VDD VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 $X=4900 $Y=1880 $D=0
M18 3 2 11 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 $X=5760 $Y=1880 $D=0
M19 5 3 VDD VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=2.4e-14 AS=1.92e-14 PD=6.2e-07 PS=5.6e-07 $X=6620 $Y=1880 $D=0
M20 VDD 4 5 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=1.92e-14 AS=2.4e-14 PD=5.6e-07 PS=6.2e-07 $X=7020 $Y=1880 $D=0
M21 17 5 3 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=2.24e-14 AS=1.92e-14 PD=6e-07 PS=5.6e-07 $X=7880 $Y=1880 $D=0
M22 VDD 1 17 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=1.92e-14 AS=2.24e-14 PD=5.6e-07 PS=6e-07 $X=8260 $Y=1880 $D=0
M23 6 1 5 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 $X=9120 $Y=1880 $D=0
M24 1 CLK_MAIN VDD VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 $X=9980 $Y=1880 $D=0
M25 2 1 VDD VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 $X=10840 $Y=1880 $D=0
M26 4 RESET VDD VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 $X=11700 $Y=1880 $D=0
M27 7 2 VDD VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=2.4e-14 AS=1.92e-14 PD=6.2e-07 PS=5.6e-07 $X=12560 $Y=1880 $D=0
M28 6 4 7 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=2.4e-14 AS=2.4e-14 PD=6.2e-07 PS=6.2e-07 $X=12960 $Y=1880 $D=0
M29 7 8 6 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=1.92e-14 AS=2.4e-14 PD=5.6e-07 PS=6.2e-07 $X=13360 $Y=1880 $D=0
M30 8 6 VDD VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 $X=14220 $Y=1880 $D=0
M31 Q 6 VDD VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 $X=15080 $Y=1880 $D=0
.ENDS
***************************************
