* SPICE NETLIST
***************************************

.SUBCKT d_flip_flop
** N=19 EP=0 IP=0 FDC=32
M0 8 7 12 12 NMOS_VTL L=5e-08 W=1e-07 AD=1.2e-14 AS=1.2e-14 PD=4.4e-07 PS=4.4e-07 $X=4040 $Y=980 $D=1
M1 9 8 12 12 NMOS_VTL L=5e-08 W=1e-07 AD=1.2e-14 AS=1.2e-14 PD=4.4e-07 PS=4.4e-07 $X=4900 $Y=980 $D=1
M2 2 1 9 12 NMOS_VTL L=5e-08 W=1e-07 AD=1.2e-14 AS=1.2e-14 PD=4.4e-07 PS=4.4e-07 $X=5760 $Y=980 $D=1
M3 16 2 12 12 NMOS_VTL L=5e-08 W=1e-07 AD=1.5e-14 AS=1.2e-14 PD=5e-07 PS=4.4e-07 $X=6620 $Y=980 $D=1
M4 3 1 16 12 NMOS_VTL L=5e-08 W=1e-07 AD=1.2e-14 AS=1.5e-14 PD=4.4e-07 PS=5e-07 $X=7020 $Y=980 $D=1
M5 17 3 2 12 NMOS_VTL L=5e-08 W=1e-07 AD=1.4e-14 AS=1.2e-14 PD=4.8e-07 PS=4.4e-07 $X=7880 $Y=980 $D=1
M6 12 1 17 12 NMOS_VTL L=5e-08 W=1e-07 AD=1.2e-14 AS=1.4e-14 PD=4.4e-07 PS=4.8e-07 $X=8260 $Y=980 $D=1
M7 4 1 3 12 NMOS_VTL L=5e-08 W=1e-07 AD=1.2e-14 AS=1.2e-14 PD=4.4e-07 PS=4.4e-07 $X=9120 $Y=980 $D=1
M8 1 10 12 12 NMOS_VTL L=5e-08 W=1e-07 AD=1.2e-14 AS=1.2e-14 PD=4.4e-07 PS=4.4e-07 $X=9980 $Y=980 $D=1
M9 1 1 12 12 NMOS_VTL L=5e-08 W=1e-07 AD=1.2e-14 AS=1.2e-14 PD=4.4e-07 PS=4.4e-07 $X=10840 $Y=980 $D=1
M10 1 11 12 12 NMOS_VTL L=5e-08 W=1e-07 AD=1.2e-14 AS=1.2e-14 PD=4.4e-07 PS=4.4e-07 $X=11700 $Y=980 $D=1
M11 18 1 12 12 NMOS_VTL L=5e-08 W=1e-07 AD=1.4e-14 AS=1.2e-14 PD=4.8e-07 PS=4.4e-07 $X=12580 $Y=980 $D=1
M12 19 1 18 12 NMOS_VTL L=5e-08 W=1e-07 AD=1.5e-14 AS=1.4e-14 PD=5e-07 PS=4.8e-07 $X=12960 $Y=980 $D=1
M13 4 6 19 12 NMOS_VTL L=5e-08 W=1e-07 AD=1.2e-14 AS=1.5e-14 PD=4.4e-07 PS=5e-07 $X=13360 $Y=980 $D=1
M14 6 4 12 12 NMOS_VTL L=5e-08 W=1e-07 AD=1.2e-14 AS=1.2e-14 PD=4.4e-07 PS=4.4e-07 $X=14220 $Y=980 $D=1
M15 14 4 12 12 NMOS_VTL L=5e-08 W=1e-07 AD=1.2e-14 AS=1.2e-14 PD=4.4e-07 PS=4.4e-07 $X=15080 $Y=980 $D=1
M16 8 7 13 13 PMOS_VTL L=5e-08 W=1.6e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 $X=4040 $Y=1880 $D=0
M17 9 8 13 13 PMOS_VTL L=5e-08 W=1.6e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 $X=4900 $Y=1880 $D=0
M18 2 1 9 13 PMOS_VTL L=5e-08 W=1.6e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 $X=5760 $Y=1880 $D=0
M19 3 2 13 13 PMOS_VTL L=5e-08 W=1.6e-07 AD=2.4e-14 AS=1.92e-14 PD=6.2e-07 PS=5.6e-07 $X=6620 $Y=1880 $D=0
M20 13 1 3 13 PMOS_VTL L=5e-08 W=1.6e-07 AD=1.92e-14 AS=2.4e-14 PD=5.6e-07 PS=6.2e-07 $X=7020 $Y=1880 $D=0
M21 15 3 2 13 PMOS_VTL L=5e-08 W=1.6e-07 AD=2.24e-14 AS=1.92e-14 PD=6e-07 PS=5.6e-07 $X=7880 $Y=1880 $D=0
M22 13 1 15 13 PMOS_VTL L=5e-08 W=1.6e-07 AD=1.92e-14 AS=2.24e-14 PD=5.6e-07 PS=6e-07 $X=8260 $Y=1880 $D=0
M23 4 1 3 13 PMOS_VTL L=5e-08 W=1.6e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 $X=9120 $Y=1880 $D=0
M24 1 10 13 13 PMOS_VTL L=5e-08 W=1.6e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 $X=9980 $Y=1880 $D=0
M25 1 1 13 13 PMOS_VTL L=5e-08 W=1.6e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 $X=10840 $Y=1880 $D=0
M26 1 11 13 13 PMOS_VTL L=5e-08 W=1.6e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 $X=11700 $Y=1880 $D=0
M27 5 1 13 13 PMOS_VTL L=5e-08 W=1.6e-07 AD=2.4e-14 AS=1.92e-14 PD=6.2e-07 PS=5.6e-07 $X=12560 $Y=1880 $D=0
M28 4 1 5 13 PMOS_VTL L=5e-08 W=1.6e-07 AD=2.4e-14 AS=2.4e-14 PD=6.2e-07 PS=6.2e-07 $X=12960 $Y=1880 $D=0
M29 5 6 4 13 PMOS_VTL L=5e-08 W=1.6e-07 AD=1.92e-14 AS=2.4e-14 PD=5.6e-07 PS=6.2e-07 $X=13360 $Y=1880 $D=0
M30 6 4 13 13 PMOS_VTL L=5e-08 W=1.6e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 $X=14220 $Y=1880 $D=0
M31 14 4 13 13 PMOS_VTL L=5e-08 W=1.6e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 $X=15080 $Y=1880 $D=0
.ENDS
***************************************
