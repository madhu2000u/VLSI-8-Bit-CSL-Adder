* SPICE NETLIST
***************************************

.SUBCKT 8_Bit_CSL_Adder VDD GND RESET S0 A0 B0 S1 A1 B1 S2 A2 B2 S3 A3 B3 S4 A4 B4 S5 A5
+ B5 S6 A6 B6 S7 A7 B7
** N=657 EP=27 IP=0 FDC=1276
M0 GND 5 S0 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.2e-14 AS=1.2e-14 PD=4.4e-07 PS=4.4e-07 $X=49850 $Y=49225 $D=1
M1 GND 10 249 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.2e-14 AS=1.2e-14 PD=4.4e-07 PS=4.4e-07 $X=50450 $Y=62980 $D=1
M2 GND 10 9 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.2e-14 AS=1.2e-14 PD=4.4e-07 PS=4.4e-07 $X=50450 $Y=63840 $D=1
M3 510 9 10 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.5e-14 AS=1.2e-14 PD=5e-07 PS=4.4e-07 $X=50450 $Y=64700 $D=1
M4 511 7 510 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.4e-14 AS=1.5e-14 PD=4.8e-07 PS=5e-07 $X=50450 $Y=65100 $D=1
M5 GND 4 511 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.2e-14 AS=1.4e-14 PD=4.4e-07 PS=4.8e-07 $X=50450 $Y=65480 $D=1
M6 GND RESET 7 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.2e-14 AS=1.2e-14 PD=4.4e-07 PS=4.4e-07 $X=50450 $Y=66360 $D=1
M7 GND 4 3 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.2e-14 AS=1.2e-14 PD=4.4e-07 PS=4.4e-07 $X=50450 $Y=67220 $D=1
M8 GND 18 4 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.2e-14 AS=1.2e-14 PD=4.4e-07 PS=4.4e-07 $X=50450 $Y=68080 $D=1
M9 11 3 10 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.2e-14 AS=1.2e-14 PD=4.4e-07 PS=4.4e-07 $X=50450 $Y=68940 $D=1
M10 512 3 GND GND NMOS_VTL L=5e-08 W=1e-07 AD=1.4e-14 AS=1.2e-14 PD=4.8e-07 PS=4.4e-07 $X=50450 $Y=69800 $D=1
M11 8 11 512 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.2e-14 AS=1.4e-14 PD=4.4e-07 PS=4.8e-07 $X=50450 $Y=70180 $D=1
M12 513 7 11 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.5e-14 AS=1.2e-14 PD=5e-07 PS=4.4e-07 $X=50450 $Y=71040 $D=1
M13 GND 8 513 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.2e-14 AS=1.5e-14 PD=4.4e-07 PS=5e-07 $X=50450 $Y=71440 $D=1
M14 250 4 8 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.2e-14 AS=1.2e-14 PD=4.4e-07 PS=4.4e-07 $X=50450 $Y=72300 $D=1
M15 GND 251 250 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.2e-14 AS=1.2e-14 PD=4.4e-07 PS=4.4e-07 $X=50450 $Y=73160 $D=1
M16 GND A0 251 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.2e-14 AS=1.2e-14 PD=4.4e-07 PS=4.4e-07 $X=50450 $Y=74020 $D=1
M17 GND 5 6 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.2e-14 AS=1.2e-14 PD=4.4e-07 PS=4.4e-07 $X=50710 $Y=49225 $D=1
M18 GND 249 253 GND NMOS_VTL L=5e-08 W=1.15e-07 AD=1.61e-14 AS=1.3225e-14 PD=5.1e-07 PS=4.6e-07 $X=50990 $Y=54715 $D=1
M19 GND 249 255 GND NMOS_VTL L=5e-08 W=1.15e-07 AD=1.61e-14 AS=1.3225e-14 PD=5.1e-07 PS=4.6e-07 $X=50990 $Y=57635 $D=1
M20 253 252 GND GND NMOS_VTL L=5e-08 W=1.15e-07 AD=1.61e-14 AS=1.61e-14 PD=5.1e-07 PS=5.1e-07 $X=51370 $Y=54715 $D=1
M21 255 252 GND GND NMOS_VTL L=5e-08 W=1.15e-07 AD=1.61e-14 AS=1.61e-14 PD=5.1e-07 PS=5.1e-07 $X=51370 $Y=57635 $D=1
M22 514 6 5 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.5e-14 AS=1.2e-14 PD=5e-07 PS=4.4e-07 $X=51570 $Y=49225 $D=1
M23 19 VDD 253 GND NMOS_VTL L=5e-08 W=1.15e-07 AD=1.61e-14 AS=1.61e-14 PD=5.1e-07 PS=5.1e-07 $X=51750 $Y=54715 $D=1
M24 20 GND 255 GND NMOS_VTL L=5e-08 W=1.15e-07 AD=1.61e-14 AS=1.61e-14 PD=5.1e-07 PS=5.1e-07 $X=51750 $Y=57635 $D=1
M25 515 17 514 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.4e-14 AS=1.5e-14 PD=4.8e-07 PS=5e-07 $X=51970 $Y=49225 $D=1
M26 516 249 19 GND NMOS_VTL L=5e-08 W=1.15e-07 AD=1.61e-14 AS=1.61e-14 PD=5.1e-07 PS=5.1e-07 $X=52130 $Y=54715 $D=1
M27 517 249 20 GND NMOS_VTL L=5e-08 W=1.15e-07 AD=1.61e-14 AS=1.61e-14 PD=5.1e-07 PS=5.1e-07 $X=52130 $Y=57635 $D=1
M28 GND 14 515 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.2e-14 AS=1.4e-14 PD=4.4e-07 PS=4.8e-07 $X=52350 $Y=49225 $D=1
M29 GND 252 516 GND NMOS_VTL L=5e-08 W=1.15e-07 AD=1.3225e-14 AS=1.61e-14 PD=4.6e-07 PS=5.1e-07 $X=52510 $Y=54715 $D=1
M30 GND 252 517 GND NMOS_VTL L=5e-08 W=1.15e-07 AD=1.3225e-14 AS=1.61e-14 PD=4.6e-07 PS=5.1e-07 $X=52510 $Y=57635 $D=1
M31 GND RESET 17 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.2e-14 AS=1.2e-14 PD=4.4e-07 PS=4.4e-07 $X=53230 $Y=49225 $D=1
M32 258 249 GND GND NMOS_VTL L=5e-08 W=1e-07 AD=1.4e-14 AS=1.15e-14 PD=4.8e-07 PS=4.3e-07 $X=53230 $Y=54745 $D=1
M33 260 249 GND GND NMOS_VTL L=5e-08 W=1e-07 AD=1.4e-14 AS=1.15e-14 PD=4.8e-07 PS=4.3e-07 $X=53230 $Y=57665 $D=1
M34 GND 252 258 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.4e-14 AS=1.4e-14 PD=4.8e-07 PS=4.8e-07 $X=53610 $Y=54745 $D=1
M35 GND 252 260 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.4e-14 AS=1.4e-14 PD=4.8e-07 PS=4.8e-07 $X=53610 $Y=57665 $D=1
M36 258 VDD GND GND NMOS_VTL L=5e-08 W=1e-07 AD=1.15e-14 AS=1.4e-14 PD=4.3e-07 PS=4.8e-07 $X=53990 $Y=54745 $D=1
M37 260 GND GND GND NMOS_VTL L=5e-08 W=1e-07 AD=1.15e-14 AS=1.4e-14 PD=4.3e-07 PS=4.8e-07 $X=53990 $Y=57665 $D=1
M38 GND 14 15 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.2e-14 AS=1.2e-14 PD=4.4e-07 PS=4.4e-07 $X=54090 $Y=49225 $D=1
M39 262 19 258 GND NMOS_VTL L=5e-08 W=9e-08 AD=1.08e-14 AS=1.125e-14 PD=4.2e-07 PS=4.3e-07 $X=54730 $Y=54745 $D=1
M40 263 20 260 GND NMOS_VTL L=5e-08 W=9e-08 AD=1.08e-14 AS=1.125e-14 PD=4.2e-07 PS=4.3e-07 $X=54730 $Y=57665 $D=1
M41 GND 18 14 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.2e-14 AS=1.2e-14 PD=4.4e-07 PS=4.4e-07 $X=54950 $Y=49225 $D=1
M42 518 VDD 262 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.4e-14 AS=1.15e-14 PD=4.8e-07 PS=4.3e-07 $X=55460 $Y=54745 $D=1
M43 519 GND 263 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.4e-14 AS=1.15e-14 PD=4.8e-07 PS=4.3e-07 $X=55460 $Y=57665 $D=1
M44 23 15 5 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.2e-14 AS=1.2e-14 PD=4.4e-07 PS=4.4e-07 $X=55810 $Y=49225 $D=1
M45 520 249 518 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.4e-14 AS=1.4e-14 PD=4.8e-07 PS=4.8e-07 $X=55840 $Y=54745 $D=1
M46 521 249 519 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.4e-14 AS=1.4e-14 PD=4.8e-07 PS=4.8e-07 $X=55840 $Y=57665 $D=1
M47 GND 27 252 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.2e-14 AS=1.2e-14 PD=4.4e-07 PS=4.4e-07 $X=55950 $Y=62980 $D=1
M48 GND 27 26 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.2e-14 AS=1.2e-14 PD=4.4e-07 PS=4.4e-07 $X=55950 $Y=63840 $D=1
M49 522 26 27 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.5e-14 AS=1.2e-14 PD=5e-07 PS=4.4e-07 $X=55950 $Y=64700 $D=1
M50 523 24 522 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.4e-14 AS=1.5e-14 PD=4.8e-07 PS=5e-07 $X=55950 $Y=65100 $D=1
M51 GND 22 523 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.2e-14 AS=1.4e-14 PD=4.4e-07 PS=4.8e-07 $X=55950 $Y=65480 $D=1
M52 GND RESET 24 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.2e-14 AS=1.2e-14 PD=4.4e-07 PS=4.4e-07 $X=55950 $Y=66360 $D=1
M53 GND 22 21 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.2e-14 AS=1.2e-14 PD=4.4e-07 PS=4.4e-07 $X=55950 $Y=67220 $D=1
M54 GND 18 22 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.2e-14 AS=1.2e-14 PD=4.4e-07 PS=4.4e-07 $X=55950 $Y=68080 $D=1
M55 28 21 27 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.2e-14 AS=1.2e-14 PD=4.4e-07 PS=4.4e-07 $X=55950 $Y=68940 $D=1
M56 524 21 GND GND NMOS_VTL L=5e-08 W=1e-07 AD=1.4e-14 AS=1.2e-14 PD=4.8e-07 PS=4.4e-07 $X=55950 $Y=69800 $D=1
M57 25 28 524 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.2e-14 AS=1.4e-14 PD=4.4e-07 PS=4.8e-07 $X=55950 $Y=70180 $D=1
M58 525 24 28 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.5e-14 AS=1.2e-14 PD=5e-07 PS=4.4e-07 $X=55950 $Y=71040 $D=1
M59 GND 25 525 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.2e-14 AS=1.5e-14 PD=4.4e-07 PS=5e-07 $X=55950 $Y=71440 $D=1
M60 264 22 25 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.2e-14 AS=1.2e-14 PD=4.4e-07 PS=4.4e-07 $X=55950 $Y=72300 $D=1
M61 GND 265 264 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.2e-14 AS=1.2e-14 PD=4.4e-07 PS=4.4e-07 $X=55950 $Y=73160 $D=1
M62 GND B0 265 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.2e-14 AS=1.2e-14 PD=4.4e-07 PS=4.4e-07 $X=55950 $Y=74020 $D=1
M63 GND 252 520 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.15e-14 AS=1.4e-14 PD=4.3e-07 PS=4.8e-07 $X=56220 $Y=54745 $D=1
M64 GND 252 521 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.15e-14 AS=1.4e-14 PD=4.3e-07 PS=4.8e-07 $X=56220 $Y=57665 $D=1
M65 526 15 GND GND NMOS_VTL L=5e-08 W=1e-07 AD=1.4e-14 AS=1.2e-14 PD=4.8e-07 PS=4.4e-07 $X=56670 $Y=49225 $D=1
M66 30 23 526 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.2e-14 AS=1.4e-14 PD=4.4e-07 PS=4.8e-07 $X=57050 $Y=49225 $D=1
M67 33 262 GND GND NMOS_VTL L=5e-08 W=1e-07 AD=1.2e-14 AS=1.2e-14 PD=4.4e-07 PS=4.4e-07 $X=57325 $Y=55295 $D=1
M68 267 GND GND GND NMOS_VTL L=5e-08 W=1e-07 AD=1.35e-14 AS=1.15e-14 PD=4.7e-07 PS=4.3e-07 $X=57350 $Y=57305 $D=1
M69 527 17 23 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.5e-14 AS=1.2e-14 PD=5e-07 PS=4.4e-07 $X=57910 $Y=49225 $D=1
M70 32 267 31 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.4e-14 AS=1.2e-14 PD=4.8e-07 PS=4.4e-07 $X=58120 $Y=57305 $D=1
M71 GND 30 527 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.2e-14 AS=1.5e-14 PD=4.4e-07 PS=5e-07 $X=58310 $Y=49225 $D=1
M72 GND 263 31 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.2e-14 AS=1.2e-14 PD=4.4e-07 PS=4.4e-07 $X=58330 $Y=58455 $D=1
M73 33 GND 32 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.15e-14 AS=1.4e-14 PD=4.3e-07 PS=4.8e-07 $X=58500 $Y=57305 $D=1
M74 268 14 30 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.2e-14 AS=1.2e-14 PD=4.4e-07 PS=4.4e-07 $X=59170 $Y=49225 $D=1
M75 GND 269 268 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.2e-14 AS=1.2e-14 PD=4.4e-07 PS=4.4e-07 $X=60030 $Y=49225 $D=1
M76 GND 32 269 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.2e-14 AS=1.2e-14 PD=4.4e-07 PS=4.4e-07 $X=60890 $Y=49225 $D=1
M77 GND 36 S1 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.2e-14 AS=1.2e-14 PD=4.4e-07 PS=4.4e-07 $X=62115 $Y=49225 $D=1
M78 GND 272 VDD GND NMOS_VTL L=5e-08 W=1e-07 AD=1.2e-14 AS=1.2e-14 PD=4.4e-07 PS=4.4e-07 $X=62155 $Y=61790 $D=1
M79 GND 41 272 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.2e-14 AS=1.2e-14 PD=4.4e-07 PS=4.4e-07 $X=62155 $Y=62975 $D=1
M80 GND 41 40 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.2e-14 AS=1.2e-14 PD=4.4e-07 PS=4.4e-07 $X=62155 $Y=63835 $D=1
M81 528 40 41 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.5e-14 AS=1.2e-14 PD=5e-07 PS=4.4e-07 $X=62155 $Y=64695 $D=1
M82 529 37 528 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.4e-14 AS=1.5e-14 PD=4.8e-07 PS=5e-07 $X=62155 $Y=65095 $D=1
M83 GND 35 529 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.2e-14 AS=1.4e-14 PD=4.4e-07 PS=4.8e-07 $X=62155 $Y=65475 $D=1
M84 GND RESET 37 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.2e-14 AS=1.2e-14 PD=4.4e-07 PS=4.4e-07 $X=62155 $Y=66355 $D=1
M85 GND 35 34 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.2e-14 AS=1.2e-14 PD=4.4e-07 PS=4.4e-07 $X=62155 $Y=67215 $D=1
M86 GND 18 35 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.2e-14 AS=1.2e-14 PD=4.4e-07 PS=4.4e-07 $X=62155 $Y=68075 $D=1
M87 42 34 41 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.2e-14 AS=1.2e-14 PD=4.4e-07 PS=4.4e-07 $X=62155 $Y=68935 $D=1
M88 530 34 GND GND NMOS_VTL L=5e-08 W=1e-07 AD=1.4e-14 AS=1.2e-14 PD=4.8e-07 PS=4.4e-07 $X=62155 $Y=69795 $D=1
M89 38 42 530 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.2e-14 AS=1.4e-14 PD=4.4e-07 PS=4.8e-07 $X=62155 $Y=70175 $D=1
M90 531 37 42 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.5e-14 AS=1.2e-14 PD=5e-07 PS=4.4e-07 $X=62155 $Y=71035 $D=1
M91 GND 38 531 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.2e-14 AS=1.5e-14 PD=4.4e-07 PS=5e-07 $X=62155 $Y=71435 $D=1
M92 273 35 38 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.2e-14 AS=1.2e-14 PD=4.4e-07 PS=4.4e-07 $X=62155 $Y=72295 $D=1
M93 GND 274 273 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.2e-14 AS=1.2e-14 PD=4.4e-07 PS=4.4e-07 $X=62155 $Y=73155 $D=1
M94 GND A1 274 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.2e-14 AS=1.2e-14 PD=4.4e-07 PS=4.4e-07 $X=62155 $Y=74015 $D=1
M95 GND VDD 276 GND NMOS_VTL L=5e-08 W=1.15e-07 AD=1.61e-14 AS=1.3225e-14 PD=5.1e-07 PS=4.6e-07 $X=62790 $Y=54715 $D=1
M96 GND VDD 278 GND NMOS_VTL L=5e-08 W=1.15e-07 AD=1.61e-14 AS=1.3225e-14 PD=5.1e-07 PS=4.6e-07 $X=62790 $Y=57795 $D=1
M97 GND 36 39 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.2e-14 AS=1.2e-14 PD=4.4e-07 PS=4.4e-07 $X=62975 $Y=49225 $D=1
M98 276 275 GND GND NMOS_VTL L=5e-08 W=1.15e-07 AD=1.61e-14 AS=1.61e-14 PD=5.1e-07 PS=5.1e-07 $X=63170 $Y=54715 $D=1
M99 278 275 GND GND NMOS_VTL L=5e-08 W=1.15e-07 AD=1.61e-14 AS=1.61e-14 PD=5.1e-07 PS=5.1e-07 $X=63170 $Y=57795 $D=1
M100 48 19 276 GND NMOS_VTL L=5e-08 W=1.15e-07 AD=1.61e-14 AS=1.61e-14 PD=5.1e-07 PS=5.1e-07 $X=63550 $Y=54715 $D=1
M101 49 20 278 GND NMOS_VTL L=5e-08 W=1.15e-07 AD=1.61e-14 AS=1.61e-14 PD=5.1e-07 PS=5.1e-07 $X=63550 $Y=57795 $D=1
M102 532 39 36 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.5e-14 AS=1.2e-14 PD=5e-07 PS=4.4e-07 $X=63835 $Y=49225 $D=1
M103 533 VDD 48 GND NMOS_VTL L=5e-08 W=1.15e-07 AD=1.61e-14 AS=1.61e-14 PD=5.1e-07 PS=5.1e-07 $X=63930 $Y=54715 $D=1
M104 534 VDD 49 GND NMOS_VTL L=5e-08 W=1.15e-07 AD=1.61e-14 AS=1.61e-14 PD=5.1e-07 PS=5.1e-07 $X=63930 $Y=57795 $D=1
M105 535 47 532 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.4e-14 AS=1.5e-14 PD=4.8e-07 PS=5e-07 $X=64235 $Y=49225 $D=1
M106 GND 275 533 GND NMOS_VTL L=5e-08 W=1.15e-07 AD=1.3225e-14 AS=1.61e-14 PD=4.6e-07 PS=5.1e-07 $X=64310 $Y=54715 $D=1
M107 GND 275 534 GND NMOS_VTL L=5e-08 W=1.15e-07 AD=1.3225e-14 AS=1.61e-14 PD=4.6e-07 PS=5.1e-07 $X=64310 $Y=57795 $D=1
M108 GND 45 535 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.2e-14 AS=1.4e-14 PD=4.4e-07 PS=4.8e-07 $X=64615 $Y=49225 $D=1
M109 280 VDD GND GND NMOS_VTL L=5e-08 W=1e-07 AD=1.4e-14 AS=1.15e-14 PD=4.8e-07 PS=4.3e-07 $X=65030 $Y=54745 $D=1
M110 282 VDD GND GND NMOS_VTL L=5e-08 W=1e-07 AD=1.4e-14 AS=1.15e-14 PD=4.8e-07 PS=4.3e-07 $X=65030 $Y=57825 $D=1
M111 GND 275 280 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.4e-14 AS=1.4e-14 PD=4.8e-07 PS=4.8e-07 $X=65410 $Y=54745 $D=1
M112 GND 275 282 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.4e-14 AS=1.4e-14 PD=4.8e-07 PS=4.8e-07 $X=65410 $Y=57825 $D=1
M113 GND RESET 47 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.2e-14 AS=1.2e-14 PD=4.4e-07 PS=4.4e-07 $X=65495 $Y=49225 $D=1
M114 280 19 GND GND NMOS_VTL L=5e-08 W=1e-07 AD=1.15e-14 AS=1.4e-14 PD=4.3e-07 PS=4.8e-07 $X=65790 $Y=54745 $D=1
M115 282 20 GND GND NMOS_VTL L=5e-08 W=1e-07 AD=1.15e-14 AS=1.4e-14 PD=4.3e-07 PS=4.8e-07 $X=65790 $Y=57825 $D=1
M116 GND 45 46 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.2e-14 AS=1.2e-14 PD=4.4e-07 PS=4.4e-07 $X=66355 $Y=49225 $D=1
M117 62 48 280 GND NMOS_VTL L=5e-08 W=9e-08 AD=1.08e-14 AS=1.125e-14 PD=4.2e-07 PS=4.3e-07 $X=66530 $Y=54745 $D=1
M118 60 49 282 GND NMOS_VTL L=5e-08 W=9e-08 AD=1.08e-14 AS=1.125e-14 PD=4.2e-07 PS=4.3e-07 $X=66530 $Y=57825 $D=1
M119 GND 18 45 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.2e-14 AS=1.2e-14 PD=4.4e-07 PS=4.4e-07 $X=67215 $Y=49225 $D=1
M120 536 19 62 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.4e-14 AS=1.15e-14 PD=4.8e-07 PS=4.3e-07 $X=67260 $Y=54745 $D=1
M121 537 20 60 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.4e-14 AS=1.15e-14 PD=4.8e-07 PS=4.3e-07 $X=67260 $Y=57825 $D=1
M122 542 VDD 536 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.4e-14 AS=1.4e-14 PD=4.8e-07 PS=4.8e-07 $X=67640 $Y=54745 $D=1
M123 543 VDD 537 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.4e-14 AS=1.4e-14 PD=4.8e-07 PS=4.8e-07 $X=67640 $Y=57825 $D=1
M124 GND 284 275 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.2e-14 AS=1.2e-14 PD=4.4e-07 PS=4.4e-07 $X=67675 $Y=61790 $D=1
M125 GND 55 284 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.2e-14 AS=1.2e-14 PD=4.4e-07 PS=4.4e-07 $X=67675 $Y=62975 $D=1
M126 GND 55 54 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.2e-14 AS=1.2e-14 PD=4.4e-07 PS=4.4e-07 $X=67675 $Y=63835 $D=1
M127 538 54 55 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.5e-14 AS=1.2e-14 PD=5e-07 PS=4.4e-07 $X=67675 $Y=64695 $D=1
M128 539 52 538 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.4e-14 AS=1.5e-14 PD=4.8e-07 PS=5e-07 $X=67675 $Y=65095 $D=1
M129 GND 51 539 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.2e-14 AS=1.4e-14 PD=4.4e-07 PS=4.8e-07 $X=67675 $Y=65475 $D=1
M130 GND RESET 52 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.2e-14 AS=1.2e-14 PD=4.4e-07 PS=4.4e-07 $X=67675 $Y=66355 $D=1
M131 GND 51 50 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.2e-14 AS=1.2e-14 PD=4.4e-07 PS=4.4e-07 $X=67675 $Y=67215 $D=1
M132 GND 18 51 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.2e-14 AS=1.2e-14 PD=4.4e-07 PS=4.4e-07 $X=67675 $Y=68075 $D=1
M133 56 50 55 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.2e-14 AS=1.2e-14 PD=4.4e-07 PS=4.4e-07 $X=67675 $Y=68935 $D=1
M134 540 50 GND GND NMOS_VTL L=5e-08 W=1e-07 AD=1.4e-14 AS=1.2e-14 PD=4.8e-07 PS=4.4e-07 $X=67675 $Y=69795 $D=1
M135 53 56 540 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.2e-14 AS=1.4e-14 PD=4.4e-07 PS=4.8e-07 $X=67675 $Y=70175 $D=1
M136 541 52 56 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.5e-14 AS=1.2e-14 PD=5e-07 PS=4.4e-07 $X=67675 $Y=71035 $D=1
M137 GND 53 541 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.2e-14 AS=1.5e-14 PD=4.4e-07 PS=5e-07 $X=67675 $Y=71435 $D=1
M138 285 51 53 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.2e-14 AS=1.2e-14 PD=4.4e-07 PS=4.4e-07 $X=67675 $Y=72295 $D=1
M139 GND 286 285 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.2e-14 AS=1.2e-14 PD=4.4e-07 PS=4.4e-07 $X=67675 $Y=73155 $D=1
M140 GND B1 286 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.2e-14 AS=1.2e-14 PD=4.4e-07 PS=4.4e-07 $X=67675 $Y=74015 $D=1
M141 GND 275 542 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.15e-14 AS=1.4e-14 PD=4.3e-07 PS=4.8e-07 $X=68020 $Y=54745 $D=1
M142 GND 275 543 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.15e-14 AS=1.4e-14 PD=4.3e-07 PS=4.8e-07 $X=68020 $Y=57825 $D=1
M143 57 46 36 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.2e-14 AS=1.2e-14 PD=4.4e-07 PS=4.4e-07 $X=68075 $Y=49225 $D=1
M144 544 46 GND GND NMOS_VTL L=5e-08 W=1e-07 AD=1.4e-14 AS=1.2e-14 PD=4.8e-07 PS=4.4e-07 $X=68935 $Y=49225 $D=1
M145 288 GND GND GND NMOS_VTL L=5e-08 W=1e-07 AD=1.35e-14 AS=1.15e-14 PD=4.7e-07 PS=4.3e-07 $X=69150 $Y=57465 $D=1
M146 59 57 544 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.2e-14 AS=1.4e-14 PD=4.4e-07 PS=4.8e-07 $X=69315 $Y=49225 $D=1
M147 61 288 60 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.4e-14 AS=1.2e-14 PD=4.8e-07 PS=4.4e-07 $X=69920 $Y=57465 $D=1
M148 545 47 57 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.5e-14 AS=1.2e-14 PD=5e-07 PS=4.4e-07 $X=70175 $Y=49225 $D=1
M149 62 GND 61 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.15e-14 AS=1.4e-14 PD=4.3e-07 PS=4.8e-07 $X=70300 $Y=57465 $D=1
M150 GND 59 545 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.2e-14 AS=1.5e-14 PD=4.4e-07 PS=5e-07 $X=70575 $Y=49225 $D=1
M151 289 45 59 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.2e-14 AS=1.2e-14 PD=4.4e-07 PS=4.4e-07 $X=71435 $Y=49225 $D=1
M152 GND 290 289 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.2e-14 AS=1.2e-14 PD=4.4e-07 PS=4.4e-07 $X=72295 $Y=49225 $D=1
M153 GND 61 290 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.2e-14 AS=1.2e-14 PD=4.4e-07 PS=4.4e-07 $X=73155 $Y=49225 $D=1
M154 GND 69 VDD GND NMOS_VTL L=5e-08 W=1e-07 AD=1.2e-14 AS=1.2e-14 PD=4.4e-07 PS=4.4e-07 $X=74050 $Y=62980 $D=1
M155 GND 69 68 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.2e-14 AS=1.2e-14 PD=4.4e-07 PS=4.4e-07 $X=74050 $Y=63840 $D=1
M156 546 68 69 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.5e-14 AS=1.2e-14 PD=5e-07 PS=4.4e-07 $X=74050 $Y=64700 $D=1
M157 547 65 546 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.4e-14 AS=1.5e-14 PD=4.8e-07 PS=5e-07 $X=74050 $Y=65100 $D=1
M158 GND 64 547 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.2e-14 AS=1.4e-14 PD=4.4e-07 PS=4.8e-07 $X=74050 $Y=65480 $D=1
M159 GND RESET 65 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.2e-14 AS=1.2e-14 PD=4.4e-07 PS=4.4e-07 $X=74050 $Y=66360 $D=1
M160 GND 64 63 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.2e-14 AS=1.2e-14 PD=4.4e-07 PS=4.4e-07 $X=74050 $Y=67220 $D=1
M161 GND 18 64 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.2e-14 AS=1.2e-14 PD=4.4e-07 PS=4.4e-07 $X=74050 $Y=68080 $D=1
M162 70 63 69 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.2e-14 AS=1.2e-14 PD=4.4e-07 PS=4.4e-07 $X=74050 $Y=68940 $D=1
M163 548 63 GND GND NMOS_VTL L=5e-08 W=1e-07 AD=1.4e-14 AS=1.2e-14 PD=4.8e-07 PS=4.4e-07 $X=74050 $Y=69800 $D=1
M164 66 70 548 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.2e-14 AS=1.4e-14 PD=4.4e-07 PS=4.8e-07 $X=74050 $Y=70180 $D=1
M165 549 65 70 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.5e-14 AS=1.2e-14 PD=5e-07 PS=4.4e-07 $X=74050 $Y=71040 $D=1
M166 GND 66 549 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.2e-14 AS=1.5e-14 PD=4.4e-07 PS=5e-07 $X=74050 $Y=71440 $D=1
M167 293 64 66 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.2e-14 AS=1.2e-14 PD=4.4e-07 PS=4.4e-07 $X=74050 $Y=72300 $D=1
M168 GND 294 293 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.2e-14 AS=1.2e-14 PD=4.4e-07 PS=4.4e-07 $X=74050 $Y=73160 $D=1
M169 GND A2 294 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.2e-14 AS=1.2e-14 PD=4.4e-07 PS=4.4e-07 $X=74050 $Y=74020 $D=1
M170 GND 67 S2 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.2e-14 AS=1.2e-14 PD=4.4e-07 PS=4.4e-07 $X=74310 $Y=49225 $D=1
M171 GND VDD 296 GND NMOS_VTL L=5e-08 W=1.15e-07 AD=1.61e-14 AS=1.3225e-14 PD=5.1e-07 PS=4.6e-07 $X=74590 $Y=54715 $D=1
M172 GND VDD 298 GND NMOS_VTL L=5e-08 W=1.15e-07 AD=1.61e-14 AS=1.3225e-14 PD=5.1e-07 PS=4.6e-07 $X=74590 $Y=57795 $D=1
M173 296 295 GND GND NMOS_VTL L=5e-08 W=1.15e-07 AD=1.61e-14 AS=1.61e-14 PD=5.1e-07 PS=5.1e-07 $X=74970 $Y=54715 $D=1
M174 298 295 GND GND NMOS_VTL L=5e-08 W=1.15e-07 AD=1.61e-14 AS=1.61e-14 PD=5.1e-07 PS=5.1e-07 $X=74970 $Y=57795 $D=1
M175 GND 67 71 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.2e-14 AS=1.2e-14 PD=4.4e-07 PS=4.4e-07 $X=75170 $Y=49225 $D=1
M176 77 48 296 GND NMOS_VTL L=5e-08 W=1.15e-07 AD=1.61e-14 AS=1.61e-14 PD=5.1e-07 PS=5.1e-07 $X=75350 $Y=54715 $D=1
M177 78 49 298 GND NMOS_VTL L=5e-08 W=1.15e-07 AD=1.61e-14 AS=1.61e-14 PD=5.1e-07 PS=5.1e-07 $X=75350 $Y=57795 $D=1
M178 550 VDD 77 GND NMOS_VTL L=5e-08 W=1.15e-07 AD=1.61e-14 AS=1.61e-14 PD=5.1e-07 PS=5.1e-07 $X=75730 $Y=54715 $D=1
M179 551 VDD 78 GND NMOS_VTL L=5e-08 W=1.15e-07 AD=1.61e-14 AS=1.61e-14 PD=5.1e-07 PS=5.1e-07 $X=75730 $Y=57795 $D=1
M180 552 71 67 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.5e-14 AS=1.2e-14 PD=5e-07 PS=4.4e-07 $X=76030 $Y=49225 $D=1
M181 GND 295 550 GND NMOS_VTL L=5e-08 W=1.15e-07 AD=1.3225e-14 AS=1.61e-14 PD=4.6e-07 PS=5.1e-07 $X=76110 $Y=54715 $D=1
M182 GND 295 551 GND NMOS_VTL L=5e-08 W=1.15e-07 AD=1.3225e-14 AS=1.61e-14 PD=4.6e-07 PS=5.1e-07 $X=76110 $Y=57795 $D=1
M183 553 76 552 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.4e-14 AS=1.5e-14 PD=4.8e-07 PS=5e-07 $X=76430 $Y=49225 $D=1
M184 GND 74 553 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.2e-14 AS=1.4e-14 PD=4.4e-07 PS=4.8e-07 $X=76810 $Y=49225 $D=1
M185 301 VDD GND GND NMOS_VTL L=5e-08 W=1e-07 AD=1.4e-14 AS=1.15e-14 PD=4.8e-07 PS=4.3e-07 $X=76830 $Y=54745 $D=1
M186 303 VDD GND GND NMOS_VTL L=5e-08 W=1e-07 AD=1.4e-14 AS=1.15e-14 PD=4.8e-07 PS=4.3e-07 $X=76830 $Y=57825 $D=1
M187 GND 295 301 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.4e-14 AS=1.4e-14 PD=4.8e-07 PS=4.8e-07 $X=77210 $Y=54745 $D=1
M188 GND 295 303 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.4e-14 AS=1.4e-14 PD=4.8e-07 PS=4.8e-07 $X=77210 $Y=57825 $D=1
M189 301 48 GND GND NMOS_VTL L=5e-08 W=1e-07 AD=1.15e-14 AS=1.4e-14 PD=4.3e-07 PS=4.8e-07 $X=77590 $Y=54745 $D=1
M190 303 49 GND GND NMOS_VTL L=5e-08 W=1e-07 AD=1.15e-14 AS=1.4e-14 PD=4.3e-07 PS=4.8e-07 $X=77590 $Y=57825 $D=1
M191 GND RESET 76 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.2e-14 AS=1.2e-14 PD=4.4e-07 PS=4.4e-07 $X=77690 $Y=49225 $D=1
M192 305 77 301 GND NMOS_VTL L=5e-08 W=9e-08 AD=1.08e-14 AS=1.125e-14 PD=4.2e-07 PS=4.3e-07 $X=78330 $Y=54745 $D=1
M193 306 78 303 GND NMOS_VTL L=5e-08 W=9e-08 AD=1.08e-14 AS=1.125e-14 PD=4.2e-07 PS=4.3e-07 $X=78330 $Y=57825 $D=1
M194 GND 74 75 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.2e-14 AS=1.2e-14 PD=4.4e-07 PS=4.4e-07 $X=78550 $Y=49225 $D=1
M195 554 48 305 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.4e-14 AS=1.15e-14 PD=4.8e-07 PS=4.3e-07 $X=79060 $Y=54745 $D=1
M196 555 49 306 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.4e-14 AS=1.15e-14 PD=4.8e-07 PS=4.3e-07 $X=79060 $Y=57825 $D=1
M197 GND 18 74 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.2e-14 AS=1.2e-14 PD=4.4e-07 PS=4.4e-07 $X=79410 $Y=49225 $D=1
M198 556 VDD 554 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.4e-14 AS=1.4e-14 PD=4.8e-07 PS=4.8e-07 $X=79440 $Y=54745 $D=1
M199 557 VDD 555 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.4e-14 AS=1.4e-14 PD=4.8e-07 PS=4.8e-07 $X=79440 $Y=57825 $D=1
M200 GND 84 295 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.2e-14 AS=1.2e-14 PD=4.4e-07 PS=4.4e-07 $X=79550 $Y=62980 $D=1
M201 GND 84 83 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.2e-14 AS=1.2e-14 PD=4.4e-07 PS=4.4e-07 $X=79550 $Y=63840 $D=1
M202 558 83 84 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.5e-14 AS=1.2e-14 PD=5e-07 PS=4.4e-07 $X=79550 $Y=64700 $D=1
M203 559 81 558 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.4e-14 AS=1.5e-14 PD=4.8e-07 PS=5e-07 $X=79550 $Y=65100 $D=1
M204 GND 80 559 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.2e-14 AS=1.4e-14 PD=4.4e-07 PS=4.8e-07 $X=79550 $Y=65480 $D=1
M205 GND RESET 81 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.2e-14 AS=1.2e-14 PD=4.4e-07 PS=4.4e-07 $X=79550 $Y=66360 $D=1
M206 GND 80 79 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.2e-14 AS=1.2e-14 PD=4.4e-07 PS=4.4e-07 $X=79550 $Y=67220 $D=1
M207 GND 18 80 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.2e-14 AS=1.2e-14 PD=4.4e-07 PS=4.4e-07 $X=79550 $Y=68080 $D=1
M208 85 79 84 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.2e-14 AS=1.2e-14 PD=4.4e-07 PS=4.4e-07 $X=79550 $Y=68940 $D=1
M209 560 79 GND GND NMOS_VTL L=5e-08 W=1e-07 AD=1.4e-14 AS=1.2e-14 PD=4.8e-07 PS=4.4e-07 $X=79550 $Y=69800 $D=1
M210 82 85 560 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.2e-14 AS=1.4e-14 PD=4.4e-07 PS=4.8e-07 $X=79550 $Y=70180 $D=1
M211 561 81 85 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.5e-14 AS=1.2e-14 PD=5e-07 PS=4.4e-07 $X=79550 $Y=71040 $D=1
M212 GND 82 561 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.2e-14 AS=1.5e-14 PD=4.4e-07 PS=5e-07 $X=79550 $Y=71440 $D=1
M213 307 80 82 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.2e-14 AS=1.2e-14 PD=4.4e-07 PS=4.4e-07 $X=79550 $Y=72300 $D=1
M214 GND 308 307 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.2e-14 AS=1.2e-14 PD=4.4e-07 PS=4.4e-07 $X=79550 $Y=73160 $D=1
M215 GND B2 308 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.2e-14 AS=1.2e-14 PD=4.4e-07 PS=4.4e-07 $X=79550 $Y=74020 $D=1
M216 GND 295 556 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.15e-14 AS=1.4e-14 PD=4.3e-07 PS=4.8e-07 $X=79820 $Y=54745 $D=1
M217 GND 295 557 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.15e-14 AS=1.4e-14 PD=4.3e-07 PS=4.8e-07 $X=79820 $Y=57825 $D=1
M218 86 75 67 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.2e-14 AS=1.2e-14 PD=4.4e-07 PS=4.4e-07 $X=80270 $Y=49225 $D=1
M219 91 305 GND GND NMOS_VTL L=5e-08 W=1e-07 AD=1.2e-14 AS=1.2e-14 PD=4.4e-07 PS=4.4e-07 $X=80925 $Y=55295 $D=1
M220 310 GND GND GND NMOS_VTL L=5e-08 W=1e-07 AD=1.35e-14 AS=1.15e-14 PD=4.7e-07 PS=4.3e-07 $X=80950 $Y=57465 $D=1
M221 562 75 GND GND NMOS_VTL L=5e-08 W=1e-07 AD=1.4e-14 AS=1.2e-14 PD=4.8e-07 PS=4.4e-07 $X=81130 $Y=49225 $D=1
M222 89 86 562 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.2e-14 AS=1.4e-14 PD=4.4e-07 PS=4.8e-07 $X=81510 $Y=49225 $D=1
M223 90 310 88 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.4e-14 AS=1.2e-14 PD=4.8e-07 PS=4.4e-07 $X=81720 $Y=57465 $D=1
M224 GND 306 88 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.2e-14 AS=1.2e-14 PD=4.4e-07 PS=4.4e-07 $X=81930 $Y=58615 $D=1
M225 91 GND 90 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.15e-14 AS=1.4e-14 PD=4.3e-07 PS=4.8e-07 $X=82100 $Y=57465 $D=1
M226 563 76 86 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.5e-14 AS=1.2e-14 PD=5e-07 PS=4.4e-07 $X=82370 $Y=49225 $D=1
M227 GND 89 563 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.2e-14 AS=1.5e-14 PD=4.4e-07 PS=5e-07 $X=82770 $Y=49225 $D=1
M228 311 74 89 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.2e-14 AS=1.2e-14 PD=4.4e-07 PS=4.4e-07 $X=83630 $Y=49225 $D=1
M229 GND 312 311 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.2e-14 AS=1.2e-14 PD=4.4e-07 PS=4.4e-07 $X=84490 $Y=49225 $D=1
M230 GND 90 312 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.2e-14 AS=1.2e-14 PD=4.4e-07 PS=4.4e-07 $X=85350 $Y=49225 $D=1
M231 GND 315 313 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.2e-14 AS=1.2e-14 PD=4.4e-07 PS=4.4e-07 $X=85755 $Y=61795 $D=1
M232 GND 97 315 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.2e-14 AS=1.2e-14 PD=4.4e-07 PS=4.4e-07 $X=85755 $Y=62980 $D=1
M233 GND 97 96 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.2e-14 AS=1.2e-14 PD=4.4e-07 PS=4.4e-07 $X=85755 $Y=63840 $D=1
M234 564 96 97 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.5e-14 AS=1.2e-14 PD=5e-07 PS=4.4e-07 $X=85755 $Y=64700 $D=1
M235 565 94 564 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.4e-14 AS=1.5e-14 PD=4.8e-07 PS=5e-07 $X=85755 $Y=65100 $D=1
M236 GND 93 565 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.2e-14 AS=1.4e-14 PD=4.4e-07 PS=4.8e-07 $X=85755 $Y=65480 $D=1
M237 GND RESET 94 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.2e-14 AS=1.2e-14 PD=4.4e-07 PS=4.4e-07 $X=85755 $Y=66360 $D=1
M238 GND 93 92 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.2e-14 AS=1.2e-14 PD=4.4e-07 PS=4.4e-07 $X=85755 $Y=67220 $D=1
M239 GND 18 93 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.2e-14 AS=1.2e-14 PD=4.4e-07 PS=4.4e-07 $X=85755 $Y=68080 $D=1
M240 98 92 97 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.2e-14 AS=1.2e-14 PD=4.4e-07 PS=4.4e-07 $X=85755 $Y=68940 $D=1
M241 566 92 GND GND NMOS_VTL L=5e-08 W=1e-07 AD=1.4e-14 AS=1.2e-14 PD=4.8e-07 PS=4.4e-07 $X=85755 $Y=69800 $D=1
M242 95 98 566 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.2e-14 AS=1.4e-14 PD=4.4e-07 PS=4.8e-07 $X=85755 $Y=70180 $D=1
M243 567 94 98 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.5e-14 AS=1.2e-14 PD=5e-07 PS=4.4e-07 $X=85755 $Y=71040 $D=1
M244 GND 95 567 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.2e-14 AS=1.5e-14 PD=4.4e-07 PS=5e-07 $X=85755 $Y=71440 $D=1
M245 316 93 95 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.2e-14 AS=1.2e-14 PD=4.4e-07 PS=4.4e-07 $X=85755 $Y=72300 $D=1
M246 GND 317 316 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.2e-14 AS=1.2e-14 PD=4.4e-07 PS=4.4e-07 $X=85755 $Y=73160 $D=1
M247 GND A3 317 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.2e-14 AS=1.2e-14 PD=4.4e-07 PS=4.4e-07 $X=85755 $Y=74020 $D=1
M248 GND 313 319 GND NMOS_VTL L=5e-08 W=1.15e-07 AD=1.61e-14 AS=1.3225e-14 PD=5.1e-07 PS=4.6e-07 $X=86390 $Y=54555 $D=1
M249 GND 313 321 GND NMOS_VTL L=5e-08 W=1.15e-07 AD=1.61e-14 AS=1.3225e-14 PD=5.1e-07 PS=4.6e-07 $X=86390 $Y=57635 $D=1
M250 GND 99 S3 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.2e-14 AS=1.2e-14 PD=4.4e-07 PS=4.4e-07 $X=86575 $Y=49225 $D=1
M251 319 318 GND GND NMOS_VTL L=5e-08 W=1.15e-07 AD=1.61e-14 AS=1.61e-14 PD=5.1e-07 PS=5.1e-07 $X=86770 $Y=54555 $D=1
M252 321 318 GND GND NMOS_VTL L=5e-08 W=1.15e-07 AD=1.61e-14 AS=1.61e-14 PD=5.1e-07 PS=5.1e-07 $X=86770 $Y=57635 $D=1
M253 106 77 319 GND NMOS_VTL L=5e-08 W=1.15e-07 AD=1.61e-14 AS=1.61e-14 PD=5.1e-07 PS=5.1e-07 $X=87150 $Y=54555 $D=1
M254 107 78 321 GND NMOS_VTL L=5e-08 W=1.15e-07 AD=1.61e-14 AS=1.61e-14 PD=5.1e-07 PS=5.1e-07 $X=87150 $Y=57635 $D=1
M255 GND 99 101 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.2e-14 AS=1.2e-14 PD=4.4e-07 PS=4.4e-07 $X=87435 $Y=49225 $D=1
M256 568 313 106 GND NMOS_VTL L=5e-08 W=1.15e-07 AD=1.61e-14 AS=1.61e-14 PD=5.1e-07 PS=5.1e-07 $X=87530 $Y=54555 $D=1
M257 569 313 107 GND NMOS_VTL L=5e-08 W=1.15e-07 AD=1.61e-14 AS=1.61e-14 PD=5.1e-07 PS=5.1e-07 $X=87530 $Y=57635 $D=1
M258 GND 318 568 GND NMOS_VTL L=5e-08 W=1.15e-07 AD=1.3225e-14 AS=1.61e-14 PD=4.6e-07 PS=5.1e-07 $X=87910 $Y=54555 $D=1
M259 GND 318 569 GND NMOS_VTL L=5e-08 W=1.15e-07 AD=1.3225e-14 AS=1.61e-14 PD=4.6e-07 PS=5.1e-07 $X=87910 $Y=57635 $D=1
M260 570 101 99 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.5e-14 AS=1.2e-14 PD=5e-07 PS=4.4e-07 $X=88295 $Y=49225 $D=1
M261 324 313 GND GND NMOS_VTL L=5e-08 W=1e-07 AD=1.4e-14 AS=1.15e-14 PD=4.8e-07 PS=4.3e-07 $X=88630 $Y=54585 $D=1
M262 326 313 GND GND NMOS_VTL L=5e-08 W=1e-07 AD=1.4e-14 AS=1.15e-14 PD=4.8e-07 PS=4.3e-07 $X=88630 $Y=57665 $D=1
M263 571 105 570 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.4e-14 AS=1.5e-14 PD=4.8e-07 PS=5e-07 $X=88695 $Y=49225 $D=1
M264 GND 318 324 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.4e-14 AS=1.4e-14 PD=4.8e-07 PS=4.8e-07 $X=89010 $Y=54585 $D=1
M265 GND 318 326 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.4e-14 AS=1.4e-14 PD=4.8e-07 PS=4.8e-07 $X=89010 $Y=57665 $D=1
M266 GND 103 571 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.2e-14 AS=1.4e-14 PD=4.4e-07 PS=4.8e-07 $X=89075 $Y=49225 $D=1
M267 324 77 GND GND NMOS_VTL L=5e-08 W=1e-07 AD=1.15e-14 AS=1.4e-14 PD=4.3e-07 PS=4.8e-07 $X=89390 $Y=54585 $D=1
M268 326 78 GND GND NMOS_VTL L=5e-08 W=1e-07 AD=1.15e-14 AS=1.4e-14 PD=4.3e-07 PS=4.8e-07 $X=89390 $Y=57665 $D=1
M269 GND RESET 105 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.2e-14 AS=1.2e-14 PD=4.4e-07 PS=4.4e-07 $X=89955 $Y=49225 $D=1
M270 120 106 324 GND NMOS_VTL L=5e-08 W=9e-08 AD=1.08e-14 AS=1.125e-14 PD=4.2e-07 PS=4.3e-07 $X=90130 $Y=54585 $D=1
M271 117 107 326 GND NMOS_VTL L=5e-08 W=9e-08 AD=1.08e-14 AS=1.125e-14 PD=4.2e-07 PS=4.3e-07 $X=90130 $Y=57665 $D=1
M272 GND 103 104 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.2e-14 AS=1.2e-14 PD=4.4e-07 PS=4.4e-07 $X=90815 $Y=49225 $D=1
M273 572 77 120 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.4e-14 AS=1.15e-14 PD=4.8e-07 PS=4.3e-07 $X=90860 $Y=54585 $D=1
M274 573 78 117 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.4e-14 AS=1.15e-14 PD=4.8e-07 PS=4.3e-07 $X=90860 $Y=57665 $D=1
M275 578 313 572 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.4e-14 AS=1.4e-14 PD=4.8e-07 PS=4.8e-07 $X=91240 $Y=54585 $D=1
M276 579 313 573 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.4e-14 AS=1.4e-14 PD=4.8e-07 PS=4.8e-07 $X=91240 $Y=57665 $D=1
M277 GND 328 318 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.2e-14 AS=1.2e-14 PD=4.4e-07 PS=4.4e-07 $X=91275 $Y=61795 $D=1
M278 GND 113 328 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.2e-14 AS=1.2e-14 PD=4.4e-07 PS=4.4e-07 $X=91275 $Y=62980 $D=1
M279 GND 113 112 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.2e-14 AS=1.2e-14 PD=4.4e-07 PS=4.4e-07 $X=91275 $Y=63840 $D=1
M280 574 112 113 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.5e-14 AS=1.2e-14 PD=5e-07 PS=4.4e-07 $X=91275 $Y=64700 $D=1
M281 575 110 574 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.4e-14 AS=1.5e-14 PD=4.8e-07 PS=5e-07 $X=91275 $Y=65100 $D=1
M282 GND 109 575 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.2e-14 AS=1.4e-14 PD=4.4e-07 PS=4.8e-07 $X=91275 $Y=65480 $D=1
M283 GND RESET 110 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.2e-14 AS=1.2e-14 PD=4.4e-07 PS=4.4e-07 $X=91275 $Y=66360 $D=1
M284 GND 109 108 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.2e-14 AS=1.2e-14 PD=4.4e-07 PS=4.4e-07 $X=91275 $Y=67220 $D=1
M285 GND 18 109 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.2e-14 AS=1.2e-14 PD=4.4e-07 PS=4.4e-07 $X=91275 $Y=68080 $D=1
M286 114 108 113 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.2e-14 AS=1.2e-14 PD=4.4e-07 PS=4.4e-07 $X=91275 $Y=68940 $D=1
M287 576 108 GND GND NMOS_VTL L=5e-08 W=1e-07 AD=1.4e-14 AS=1.2e-14 PD=4.8e-07 PS=4.4e-07 $X=91275 $Y=69800 $D=1
M288 111 114 576 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.2e-14 AS=1.4e-14 PD=4.4e-07 PS=4.8e-07 $X=91275 $Y=70180 $D=1
M289 577 110 114 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.5e-14 AS=1.2e-14 PD=5e-07 PS=4.4e-07 $X=91275 $Y=71040 $D=1
M290 GND 111 577 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.2e-14 AS=1.5e-14 PD=4.4e-07 PS=5e-07 $X=91275 $Y=71440 $D=1
M291 329 109 111 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.2e-14 AS=1.2e-14 PD=4.4e-07 PS=4.4e-07 $X=91275 $Y=72300 $D=1
M292 GND 330 329 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.2e-14 AS=1.2e-14 PD=4.4e-07 PS=4.4e-07 $X=91275 $Y=73160 $D=1
M293 GND B3 330 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.2e-14 AS=1.2e-14 PD=4.4e-07 PS=4.4e-07 $X=91275 $Y=74020 $D=1
M294 GND 318 578 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.15e-14 AS=1.4e-14 PD=4.3e-07 PS=4.8e-07 $X=91620 $Y=54585 $D=1
M295 GND 318 579 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.15e-14 AS=1.4e-14 PD=4.3e-07 PS=4.8e-07 $X=91620 $Y=57665 $D=1
M296 GND 18 103 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.2e-14 AS=1.2e-14 PD=4.4e-07 PS=4.4e-07 $X=91675 $Y=49225 $D=1
M297 116 104 99 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.2e-14 AS=1.2e-14 PD=4.4e-07 PS=4.4e-07 $X=92535 $Y=49225 $D=1
M298 332 GND GND GND NMOS_VTL L=5e-08 W=1e-07 AD=1.35e-14 AS=1.15e-14 PD=4.7e-07 PS=4.3e-07 $X=92750 $Y=57305 $D=1
M299 580 104 GND GND NMOS_VTL L=5e-08 W=1e-07 AD=1.4e-14 AS=1.2e-14 PD=4.8e-07 PS=4.4e-07 $X=93395 $Y=49225 $D=1
M300 118 332 117 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.4e-14 AS=1.2e-14 PD=4.8e-07 PS=4.4e-07 $X=93520 $Y=57305 $D=1
M301 119 116 580 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.2e-14 AS=1.4e-14 PD=4.4e-07 PS=4.8e-07 $X=93775 $Y=49225 $D=1
M302 120 GND 118 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.15e-14 AS=1.4e-14 PD=4.3e-07 PS=4.8e-07 $X=93900 $Y=57305 $D=1
M303 581 105 116 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.5e-14 AS=1.2e-14 PD=5e-07 PS=4.4e-07 $X=94635 $Y=49225 $D=1
M304 GND 119 581 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.2e-14 AS=1.5e-14 PD=4.4e-07 PS=5e-07 $X=95035 $Y=49225 $D=1
M305 333 GND GND GND NMOS_VTL L=5e-08 W=1e-07 AD=1.35e-14 AS=1.15e-14 PD=4.7e-07 PS=4.3e-07 $X=95855 $Y=57280 $D=1
M306 334 103 119 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.2e-14 AS=1.2e-14 PD=4.4e-07 PS=4.4e-07 $X=95895 $Y=49225 $D=1
M307 121 333 107 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.4e-14 AS=1.2e-14 PD=4.8e-07 PS=4.4e-07 $X=96625 $Y=57280 $D=1
M308 GND 335 334 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.2e-14 AS=1.2e-14 PD=4.4e-07 PS=4.4e-07 $X=96755 $Y=49225 $D=1
M309 106 GND 121 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.15e-14 AS=1.4e-14 PD=4.3e-07 PS=4.8e-07 $X=97005 $Y=57280 $D=1
M310 GND 118 335 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.2e-14 AS=1.2e-14 PD=4.4e-07 PS=4.4e-07 $X=97615 $Y=49225 $D=1
M311 GND 122 S4 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.2e-14 AS=1.2e-14 PD=4.4e-07 PS=4.4e-07 $X=99550 $Y=49225 $D=1
M312 GND 122 123 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.2e-14 AS=1.2e-14 PD=4.4e-07 PS=4.4e-07 $X=100410 $Y=49225 $D=1
M313 GND 130 338 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.2e-14 AS=1.2e-14 PD=4.4e-07 PS=4.4e-07 $X=100920 $Y=62980 $D=1
M314 GND 130 129 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.2e-14 AS=1.2e-14 PD=4.4e-07 PS=4.4e-07 $X=100920 $Y=63840 $D=1
M315 582 129 130 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.5e-14 AS=1.2e-14 PD=5e-07 PS=4.4e-07 $X=100920 $Y=64700 $D=1
M316 583 127 582 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.4e-14 AS=1.5e-14 PD=4.8e-07 PS=5e-07 $X=100920 $Y=65100 $D=1
M317 GND 125 583 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.2e-14 AS=1.4e-14 PD=4.4e-07 PS=4.8e-07 $X=100920 $Y=65480 $D=1
M318 GND RESET 127 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.2e-14 AS=1.2e-14 PD=4.4e-07 PS=4.4e-07 $X=100920 $Y=66360 $D=1
M319 GND 125 124 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.2e-14 AS=1.2e-14 PD=4.4e-07 PS=4.4e-07 $X=100920 $Y=67220 $D=1
M320 GND 18 125 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.2e-14 AS=1.2e-14 PD=4.4e-07 PS=4.4e-07 $X=100920 $Y=68080 $D=1
M321 131 124 130 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.2e-14 AS=1.2e-14 PD=4.4e-07 PS=4.4e-07 $X=100920 $Y=68940 $D=1
M322 584 124 GND GND NMOS_VTL L=5e-08 W=1e-07 AD=1.4e-14 AS=1.2e-14 PD=4.8e-07 PS=4.4e-07 $X=100920 $Y=69800 $D=1
M323 128 131 584 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.2e-14 AS=1.4e-14 PD=4.4e-07 PS=4.8e-07 $X=100920 $Y=70180 $D=1
M324 585 127 131 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.5e-14 AS=1.2e-14 PD=5e-07 PS=4.4e-07 $X=100920 $Y=71040 $D=1
M325 GND 128 585 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.2e-14 AS=1.5e-14 PD=4.4e-07 PS=5e-07 $X=100920 $Y=71440 $D=1
M326 339 125 128 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.2e-14 AS=1.2e-14 PD=4.4e-07 PS=4.4e-07 $X=100920 $Y=72300 $D=1
M327 GND 340 339 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.2e-14 AS=1.2e-14 PD=4.4e-07 PS=4.4e-07 $X=100920 $Y=73160 $D=1
M328 GND A4 340 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.2e-14 AS=1.2e-14 PD=4.4e-07 PS=4.4e-07 $X=100920 $Y=74020 $D=1
M329 586 123 122 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.5e-14 AS=1.2e-14 PD=5e-07 PS=4.4e-07 $X=101270 $Y=49225 $D=1
M330 GND 338 342 GND NMOS_VTL L=5e-08 W=1.15e-07 AD=1.61e-14 AS=1.3225e-14 PD=5.1e-07 PS=4.6e-07 $X=101460 $Y=54715 $D=1
M331 GND 338 344 GND NMOS_VTL L=5e-08 W=1.15e-07 AD=1.61e-14 AS=1.3225e-14 PD=5.1e-07 PS=4.6e-07 $X=101460 $Y=57635 $D=1
M332 587 135 586 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.4e-14 AS=1.5e-14 PD=4.8e-07 PS=5e-07 $X=101670 $Y=49225 $D=1
M333 342 341 GND GND NMOS_VTL L=5e-08 W=1.15e-07 AD=1.61e-14 AS=1.61e-14 PD=5.1e-07 PS=5.1e-07 $X=101840 $Y=54715 $D=1
M334 344 341 GND GND NMOS_VTL L=5e-08 W=1.15e-07 AD=1.61e-14 AS=1.61e-14 PD=5.1e-07 PS=5.1e-07 $X=101840 $Y=57635 $D=1
M335 GND 133 587 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.2e-14 AS=1.4e-14 PD=4.4e-07 PS=4.8e-07 $X=102050 $Y=49225 $D=1
M336 136 147 342 GND NMOS_VTL L=5e-08 W=1.15e-07 AD=1.61e-14 AS=1.61e-14 PD=5.1e-07 PS=5.1e-07 $X=102220 $Y=54715 $D=1
M337 137 GND 344 GND NMOS_VTL L=5e-08 W=1.15e-07 AD=1.61e-14 AS=1.61e-14 PD=5.1e-07 PS=5.1e-07 $X=102220 $Y=57635 $D=1
M338 588 338 136 GND NMOS_VTL L=5e-08 W=1.15e-07 AD=1.61e-14 AS=1.61e-14 PD=5.1e-07 PS=5.1e-07 $X=102600 $Y=54715 $D=1
M339 589 338 137 GND NMOS_VTL L=5e-08 W=1.15e-07 AD=1.61e-14 AS=1.61e-14 PD=5.1e-07 PS=5.1e-07 $X=102600 $Y=57635 $D=1
M340 GND RESET 135 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.2e-14 AS=1.2e-14 PD=4.4e-07 PS=4.4e-07 $X=102930 $Y=49225 $D=1
M341 GND 341 588 GND NMOS_VTL L=5e-08 W=1.15e-07 AD=1.3225e-14 AS=1.61e-14 PD=4.6e-07 PS=5.1e-07 $X=102980 $Y=54715 $D=1
M342 GND 341 589 GND NMOS_VTL L=5e-08 W=1.15e-07 AD=1.3225e-14 AS=1.61e-14 PD=4.6e-07 PS=5.1e-07 $X=102980 $Y=57635 $D=1
M343 347 338 GND GND NMOS_VTL L=5e-08 W=1e-07 AD=1.4e-14 AS=1.15e-14 PD=4.8e-07 PS=4.3e-07 $X=103700 $Y=54745 $D=1
M344 349 338 GND GND NMOS_VTL L=5e-08 W=1e-07 AD=1.4e-14 AS=1.15e-14 PD=4.8e-07 PS=4.3e-07 $X=103700 $Y=57665 $D=1
M345 GND 133 134 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.2e-14 AS=1.2e-14 PD=4.4e-07 PS=4.4e-07 $X=103790 $Y=49225 $D=1
M346 GND 341 347 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.4e-14 AS=1.4e-14 PD=4.8e-07 PS=4.8e-07 $X=104080 $Y=54745 $D=1
M347 GND 341 349 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.4e-14 AS=1.4e-14 PD=4.8e-07 PS=4.8e-07 $X=104080 $Y=57665 $D=1
M348 347 147 GND GND NMOS_VTL L=5e-08 W=1e-07 AD=1.15e-14 AS=1.4e-14 PD=4.3e-07 PS=4.8e-07 $X=104460 $Y=54745 $D=1
M349 349 GND GND GND NMOS_VTL L=5e-08 W=1e-07 AD=1.15e-14 AS=1.4e-14 PD=4.3e-07 PS=4.8e-07 $X=104460 $Y=57665 $D=1
M350 GND 18 133 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.2e-14 AS=1.2e-14 PD=4.4e-07 PS=4.4e-07 $X=104650 $Y=49225 $D=1
M351 351 136 347 GND NMOS_VTL L=5e-08 W=9e-08 AD=1.08e-14 AS=1.125e-14 PD=4.2e-07 PS=4.3e-07 $X=105200 $Y=54745 $D=1
M352 352 137 349 GND NMOS_VTL L=5e-08 W=9e-08 AD=1.08e-14 AS=1.125e-14 PD=4.2e-07 PS=4.3e-07 $X=105200 $Y=57665 $D=1
M353 139 134 122 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.2e-14 AS=1.2e-14 PD=4.4e-07 PS=4.4e-07 $X=105510 $Y=49225 $D=1
M354 590 147 351 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.4e-14 AS=1.15e-14 PD=4.8e-07 PS=4.3e-07 $X=105930 $Y=54745 $D=1
M355 591 GND 352 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.4e-14 AS=1.15e-14 PD=4.8e-07 PS=4.3e-07 $X=105930 $Y=57665 $D=1
M356 592 338 590 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.4e-14 AS=1.4e-14 PD=4.8e-07 PS=4.8e-07 $X=106310 $Y=54745 $D=1
M357 593 338 591 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.4e-14 AS=1.4e-14 PD=4.8e-07 PS=4.8e-07 $X=106310 $Y=57665 $D=1
M358 598 134 GND GND NMOS_VTL L=5e-08 W=1e-07 AD=1.4e-14 AS=1.2e-14 PD=4.8e-07 PS=4.4e-07 $X=106370 $Y=49225 $D=1
M359 GND 144 341 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.2e-14 AS=1.2e-14 PD=4.4e-07 PS=4.4e-07 $X=106420 $Y=62980 $D=1
M360 GND 144 143 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.2e-14 AS=1.2e-14 PD=4.4e-07 PS=4.4e-07 $X=106420 $Y=63840 $D=1
M361 594 143 144 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.5e-14 AS=1.2e-14 PD=5e-07 PS=4.4e-07 $X=106420 $Y=64700 $D=1
M362 595 141 594 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.4e-14 AS=1.5e-14 PD=4.8e-07 PS=5e-07 $X=106420 $Y=65100 $D=1
M363 GND 140 595 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.2e-14 AS=1.4e-14 PD=4.4e-07 PS=4.8e-07 $X=106420 $Y=65480 $D=1
M364 GND RESET 141 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.2e-14 AS=1.2e-14 PD=4.4e-07 PS=4.4e-07 $X=106420 $Y=66360 $D=1
M365 GND 140 138 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.2e-14 AS=1.2e-14 PD=4.4e-07 PS=4.4e-07 $X=106420 $Y=67220 $D=1
M366 GND 18 140 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.2e-14 AS=1.2e-14 PD=4.4e-07 PS=4.4e-07 $X=106420 $Y=68080 $D=1
M367 145 138 144 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.2e-14 AS=1.2e-14 PD=4.4e-07 PS=4.4e-07 $X=106420 $Y=68940 $D=1
M368 596 138 GND GND NMOS_VTL L=5e-08 W=1e-07 AD=1.4e-14 AS=1.2e-14 PD=4.8e-07 PS=4.4e-07 $X=106420 $Y=69800 $D=1
M369 142 145 596 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.2e-14 AS=1.4e-14 PD=4.4e-07 PS=4.8e-07 $X=106420 $Y=70180 $D=1
M370 597 141 145 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.5e-14 AS=1.2e-14 PD=5e-07 PS=4.4e-07 $X=106420 $Y=71040 $D=1
M371 GND 142 597 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.2e-14 AS=1.5e-14 PD=4.4e-07 PS=5e-07 $X=106420 $Y=71440 $D=1
M372 353 140 142 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.2e-14 AS=1.2e-14 PD=4.4e-07 PS=4.4e-07 $X=106420 $Y=72300 $D=1
M373 GND 354 353 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.2e-14 AS=1.2e-14 PD=4.4e-07 PS=4.4e-07 $X=106420 $Y=73160 $D=1
M374 GND B4 354 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.2e-14 AS=1.2e-14 PD=4.4e-07 PS=4.4e-07 $X=106420 $Y=74020 $D=1
M375 GND 341 592 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.15e-14 AS=1.4e-14 PD=4.3e-07 PS=4.8e-07 $X=106690 $Y=54745 $D=1
M376 GND 341 593 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.15e-14 AS=1.4e-14 PD=4.3e-07 PS=4.8e-07 $X=106690 $Y=57665 $D=1
M377 146 139 598 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.2e-14 AS=1.4e-14 PD=4.4e-07 PS=4.8e-07 $X=106750 $Y=49225 $D=1
M378 599 135 139 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.5e-14 AS=1.2e-14 PD=5e-07 PS=4.4e-07 $X=107610 $Y=49225 $D=1
M379 151 351 GND GND NMOS_VTL L=5e-08 W=1e-07 AD=1.2e-14 AS=1.2e-14 PD=4.4e-07 PS=4.4e-07 $X=107795 $Y=55295 $D=1
M380 356 121 GND GND NMOS_VTL L=5e-08 W=1e-07 AD=1.35e-14 AS=1.15e-14 PD=4.7e-07 PS=4.3e-07 $X=107820 $Y=57305 $D=1
M381 GND 146 599 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.2e-14 AS=1.5e-14 PD=4.4e-07 PS=5e-07 $X=108010 $Y=49225 $D=1
M382 150 356 149 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.4e-14 AS=1.2e-14 PD=4.8e-07 PS=4.4e-07 $X=108590 $Y=57305 $D=1
M383 GND 352 149 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.2e-14 AS=1.2e-14 PD=4.4e-07 PS=4.4e-07 $X=108800 $Y=58455 $D=1
M384 357 133 146 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.2e-14 AS=1.2e-14 PD=4.4e-07 PS=4.4e-07 $X=108870 $Y=49225 $D=1
M385 151 121 150 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.15e-14 AS=1.4e-14 PD=4.3e-07 PS=4.8e-07 $X=108970 $Y=57305 $D=1
M386 GND 358 357 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.2e-14 AS=1.2e-14 PD=4.4e-07 PS=4.4e-07 $X=109730 $Y=49225 $D=1
M387 GND 150 358 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.2e-14 AS=1.2e-14 PD=4.4e-07 PS=4.4e-07 $X=110590 $Y=49225 $D=1
M388 GND 154 S5 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.2e-14 AS=1.2e-14 PD=4.4e-07 PS=4.4e-07 $X=111970 $Y=49225 $D=1
M389 GND 362 361 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.2e-14 AS=1.2e-14 PD=4.4e-07 PS=4.4e-07 $X=112625 $Y=61795 $D=1
M390 GND 159 362 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.2e-14 AS=1.2e-14 PD=4.4e-07 PS=4.4e-07 $X=112625 $Y=62980 $D=1
M391 GND 159 158 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.2e-14 AS=1.2e-14 PD=4.4e-07 PS=4.4e-07 $X=112625 $Y=63840 $D=1
M392 600 158 159 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.5e-14 AS=1.2e-14 PD=5e-07 PS=4.4e-07 $X=112625 $Y=64700 $D=1
M393 601 156 600 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.4e-14 AS=1.5e-14 PD=4.8e-07 PS=5e-07 $X=112625 $Y=65100 $D=1
M394 GND 153 601 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.2e-14 AS=1.4e-14 PD=4.4e-07 PS=4.8e-07 $X=112625 $Y=65480 $D=1
M395 GND RESET 156 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.2e-14 AS=1.2e-14 PD=4.4e-07 PS=4.4e-07 $X=112625 $Y=66360 $D=1
M396 GND 153 152 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.2e-14 AS=1.2e-14 PD=4.4e-07 PS=4.4e-07 $X=112625 $Y=67220 $D=1
M397 GND 18 153 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.2e-14 AS=1.2e-14 PD=4.4e-07 PS=4.4e-07 $X=112625 $Y=68080 $D=1
M398 160 152 159 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.2e-14 AS=1.2e-14 PD=4.4e-07 PS=4.4e-07 $X=112625 $Y=68940 $D=1
M399 602 152 GND GND NMOS_VTL L=5e-08 W=1e-07 AD=1.4e-14 AS=1.2e-14 PD=4.8e-07 PS=4.4e-07 $X=112625 $Y=69800 $D=1
M400 157 160 602 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.2e-14 AS=1.4e-14 PD=4.4e-07 PS=4.8e-07 $X=112625 $Y=70180 $D=1
M401 603 156 160 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.5e-14 AS=1.2e-14 PD=5e-07 PS=4.4e-07 $X=112625 $Y=71040 $D=1
M402 GND 157 603 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.2e-14 AS=1.5e-14 PD=4.4e-07 PS=5e-07 $X=112625 $Y=71440 $D=1
M403 363 153 157 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.2e-14 AS=1.2e-14 PD=4.4e-07 PS=4.4e-07 $X=112625 $Y=72300 $D=1
M404 GND 364 363 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.2e-14 AS=1.2e-14 PD=4.4e-07 PS=4.4e-07 $X=112625 $Y=73160 $D=1
M405 GND A5 364 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.2e-14 AS=1.2e-14 PD=4.4e-07 PS=4.4e-07 $X=112625 $Y=74020 $D=1
M406 GND 154 155 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.2e-14 AS=1.2e-14 PD=4.4e-07 PS=4.4e-07 $X=112830 $Y=49225 $D=1
M407 GND 361 366 GND NMOS_VTL L=5e-08 W=1.15e-07 AD=1.61e-14 AS=1.3225e-14 PD=5.1e-07 PS=4.6e-07 $X=113260 $Y=54505 $D=1
M408 GND 361 368 GND NMOS_VTL L=5e-08 W=1.15e-07 AD=1.61e-14 AS=1.3225e-14 PD=5.1e-07 PS=4.6e-07 $X=113260 $Y=57585 $D=1
M409 366 365 GND GND NMOS_VTL L=5e-08 W=1.15e-07 AD=1.61e-14 AS=1.61e-14 PD=5.1e-07 PS=5.1e-07 $X=113640 $Y=54505 $D=1
M410 368 365 GND GND NMOS_VTL L=5e-08 W=1.15e-07 AD=1.61e-14 AS=1.61e-14 PD=5.1e-07 PS=5.1e-07 $X=113640 $Y=57585 $D=1
M411 604 155 154 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.5e-14 AS=1.2e-14 PD=5e-07 PS=4.4e-07 $X=113690 $Y=49225 $D=1
M412 166 136 366 GND NMOS_VTL L=5e-08 W=1.15e-07 AD=1.61e-14 AS=1.61e-14 PD=5.1e-07 PS=5.1e-07 $X=114020 $Y=54505 $D=1
M413 167 137 368 GND NMOS_VTL L=5e-08 W=1.15e-07 AD=1.61e-14 AS=1.61e-14 PD=5.1e-07 PS=5.1e-07 $X=114020 $Y=57585 $D=1
M414 605 165 604 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.4e-14 AS=1.5e-14 PD=4.8e-07 PS=5e-07 $X=114090 $Y=49225 $D=1
M415 606 361 166 GND NMOS_VTL L=5e-08 W=1.15e-07 AD=1.61e-14 AS=1.61e-14 PD=5.1e-07 PS=5.1e-07 $X=114400 $Y=54505 $D=1
M416 607 361 167 GND NMOS_VTL L=5e-08 W=1.15e-07 AD=1.61e-14 AS=1.61e-14 PD=5.1e-07 PS=5.1e-07 $X=114400 $Y=57585 $D=1
M417 GND 163 605 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.2e-14 AS=1.4e-14 PD=4.4e-07 PS=4.8e-07 $X=114470 $Y=49225 $D=1
M418 GND 365 606 GND NMOS_VTL L=5e-08 W=1.15e-07 AD=1.3225e-14 AS=1.61e-14 PD=4.6e-07 PS=5.1e-07 $X=114780 $Y=54505 $D=1
M419 GND 365 607 GND NMOS_VTL L=5e-08 W=1.15e-07 AD=1.3225e-14 AS=1.61e-14 PD=4.6e-07 PS=5.1e-07 $X=114780 $Y=57585 $D=1
M420 GND RESET 165 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.2e-14 AS=1.2e-14 PD=4.4e-07 PS=4.4e-07 $X=115350 $Y=49225 $D=1
M421 371 361 GND GND NMOS_VTL L=5e-08 W=1e-07 AD=1.4e-14 AS=1.15e-14 PD=4.8e-07 PS=4.3e-07 $X=115500 $Y=54535 $D=1
M422 373 361 GND GND NMOS_VTL L=5e-08 W=1e-07 AD=1.4e-14 AS=1.15e-14 PD=4.8e-07 PS=4.3e-07 $X=115500 $Y=57615 $D=1
M423 GND 365 371 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.4e-14 AS=1.4e-14 PD=4.8e-07 PS=4.8e-07 $X=115880 $Y=54535 $D=1
M424 GND 365 373 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.4e-14 AS=1.4e-14 PD=4.8e-07 PS=4.8e-07 $X=115880 $Y=57615 $D=1
M425 GND 163 164 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.2e-14 AS=1.2e-14 PD=4.4e-07 PS=4.4e-07 $X=116210 $Y=49225 $D=1
M426 371 136 GND GND NMOS_VTL L=5e-08 W=1e-07 AD=1.15e-14 AS=1.4e-14 PD=4.3e-07 PS=4.8e-07 $X=116260 $Y=54535 $D=1
M427 373 137 GND GND NMOS_VTL L=5e-08 W=1e-07 AD=1.15e-14 AS=1.4e-14 PD=4.3e-07 PS=4.8e-07 $X=116260 $Y=57615 $D=1
M428 375 166 371 GND NMOS_VTL L=5e-08 W=9e-08 AD=1.08e-14 AS=1.125e-14 PD=4.2e-07 PS=4.3e-07 $X=117000 $Y=54535 $D=1
M429 178 167 373 GND NMOS_VTL L=5e-08 W=9e-08 AD=1.08e-14 AS=1.125e-14 PD=4.2e-07 PS=4.3e-07 $X=117000 $Y=57615 $D=1
M430 GND 18 163 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.2e-14 AS=1.2e-14 PD=4.4e-07 PS=4.4e-07 $X=117070 $Y=49225 $D=1
M431 608 136 375 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.4e-14 AS=1.15e-14 PD=4.8e-07 PS=4.3e-07 $X=117730 $Y=54535 $D=1
M432 609 137 178 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.4e-14 AS=1.15e-14 PD=4.8e-07 PS=4.3e-07 $X=117730 $Y=57615 $D=1
M433 170 164 154 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.2e-14 AS=1.2e-14 PD=4.4e-07 PS=4.4e-07 $X=117930 $Y=49225 $D=1
M434 614 361 608 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.4e-14 AS=1.4e-14 PD=4.8e-07 PS=4.8e-07 $X=118110 $Y=54535 $D=1
M435 615 361 609 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.4e-14 AS=1.4e-14 PD=4.8e-07 PS=4.8e-07 $X=118110 $Y=57615 $D=1
M436 GND 376 365 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.2e-14 AS=1.2e-14 PD=4.4e-07 PS=4.4e-07 $X=118145 $Y=61795 $D=1
M437 GND 174 376 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.2e-14 AS=1.2e-14 PD=4.4e-07 PS=4.4e-07 $X=118145 $Y=62980 $D=1
M438 GND 174 173 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.2e-14 AS=1.2e-14 PD=4.4e-07 PS=4.4e-07 $X=118145 $Y=63840 $D=1
M439 610 173 174 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.5e-14 AS=1.2e-14 PD=5e-07 PS=4.4e-07 $X=118145 $Y=64700 $D=1
M440 611 171 610 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.4e-14 AS=1.5e-14 PD=4.8e-07 PS=5e-07 $X=118145 $Y=65100 $D=1
M441 GND 169 611 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.2e-14 AS=1.4e-14 PD=4.4e-07 PS=4.8e-07 $X=118145 $Y=65480 $D=1
M442 GND RESET 171 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.2e-14 AS=1.2e-14 PD=4.4e-07 PS=4.4e-07 $X=118145 $Y=66360 $D=1
M443 GND 169 168 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.2e-14 AS=1.2e-14 PD=4.4e-07 PS=4.4e-07 $X=118145 $Y=67220 $D=1
M444 GND 18 169 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.2e-14 AS=1.2e-14 PD=4.4e-07 PS=4.4e-07 $X=118145 $Y=68080 $D=1
M445 175 168 174 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.2e-14 AS=1.2e-14 PD=4.4e-07 PS=4.4e-07 $X=118145 $Y=68940 $D=1
M446 612 168 GND GND NMOS_VTL L=5e-08 W=1e-07 AD=1.4e-14 AS=1.2e-14 PD=4.8e-07 PS=4.4e-07 $X=118145 $Y=69800 $D=1
M447 172 175 612 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.2e-14 AS=1.4e-14 PD=4.4e-07 PS=4.8e-07 $X=118145 $Y=70180 $D=1
M448 613 171 175 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.5e-14 AS=1.2e-14 PD=5e-07 PS=4.4e-07 $X=118145 $Y=71040 $D=1
M449 GND 172 613 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.2e-14 AS=1.5e-14 PD=4.4e-07 PS=5e-07 $X=118145 $Y=71440 $D=1
M450 377 169 172 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.2e-14 AS=1.2e-14 PD=4.4e-07 PS=4.4e-07 $X=118145 $Y=72300 $D=1
M451 GND 378 377 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.2e-14 AS=1.2e-14 PD=4.4e-07 PS=4.4e-07 $X=118145 $Y=73160 $D=1
M452 GND B5 378 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.2e-14 AS=1.2e-14 PD=4.4e-07 PS=4.4e-07 $X=118145 $Y=74020 $D=1
M453 GND 365 614 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.15e-14 AS=1.4e-14 PD=4.3e-07 PS=4.8e-07 $X=118490 $Y=54535 $D=1
M454 GND 365 615 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.15e-14 AS=1.4e-14 PD=4.3e-07 PS=4.8e-07 $X=118490 $Y=57615 $D=1
M455 616 164 GND GND NMOS_VTL L=5e-08 W=1e-07 AD=1.4e-14 AS=1.2e-14 PD=4.8e-07 PS=4.4e-07 $X=118790 $Y=49225 $D=1
M456 177 170 616 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.2e-14 AS=1.4e-14 PD=4.4e-07 PS=4.8e-07 $X=119170 $Y=49225 $D=1
M457 381 121 GND GND NMOS_VTL L=5e-08 W=1e-07 AD=1.35e-14 AS=1.15e-14 PD=4.7e-07 PS=4.3e-07 $X=119620 $Y=57255 $D=1
M458 617 165 170 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.5e-14 AS=1.2e-14 PD=5e-07 PS=4.4e-07 $X=120030 $Y=49225 $D=1
M459 179 381 178 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.4e-14 AS=1.2e-14 PD=4.8e-07 PS=4.4e-07 $X=120390 $Y=57255 $D=1
M460 GND 177 617 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.2e-14 AS=1.5e-14 PD=4.4e-07 PS=5e-07 $X=120430 $Y=49225 $D=1
M461 180 121 179 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.15e-14 AS=1.4e-14 PD=4.3e-07 PS=4.8e-07 $X=120770 $Y=57255 $D=1
M462 382 163 177 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.2e-14 AS=1.2e-14 PD=4.4e-07 PS=4.4e-07 $X=121290 $Y=49225 $D=1
M463 GND 383 382 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.2e-14 AS=1.2e-14 PD=4.4e-07 PS=4.4e-07 $X=122150 $Y=49225 $D=1
M464 GND 179 383 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.2e-14 AS=1.2e-14 PD=4.4e-07 PS=4.4e-07 $X=123010 $Y=49225 $D=1
M465 GND 188 386 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.2e-14 AS=1.2e-14 PD=4.4e-07 PS=4.4e-07 $X=124520 $Y=62980 $D=1
M466 GND 188 187 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.2e-14 AS=1.2e-14 PD=4.4e-07 PS=4.4e-07 $X=124520 $Y=63840 $D=1
M467 618 187 188 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.5e-14 AS=1.2e-14 PD=5e-07 PS=4.4e-07 $X=124520 $Y=64700 $D=1
M468 619 184 618 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.4e-14 AS=1.5e-14 PD=4.8e-07 PS=5e-07 $X=124520 $Y=65100 $D=1
M469 GND 182 619 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.2e-14 AS=1.4e-14 PD=4.4e-07 PS=4.8e-07 $X=124520 $Y=65480 $D=1
M470 GND RESET 184 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.2e-14 AS=1.2e-14 PD=4.4e-07 PS=4.4e-07 $X=124520 $Y=66360 $D=1
M471 GND 182 181 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.2e-14 AS=1.2e-14 PD=4.4e-07 PS=4.4e-07 $X=124520 $Y=67220 $D=1
M472 GND 18 182 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.2e-14 AS=1.2e-14 PD=4.4e-07 PS=4.4e-07 $X=124520 $Y=68080 $D=1
M473 189 181 188 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.2e-14 AS=1.2e-14 PD=4.4e-07 PS=4.4e-07 $X=124520 $Y=68940 $D=1
M474 620 181 GND GND NMOS_VTL L=5e-08 W=1e-07 AD=1.4e-14 AS=1.2e-14 PD=4.8e-07 PS=4.4e-07 $X=124520 $Y=69800 $D=1
M475 185 189 620 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.2e-14 AS=1.4e-14 PD=4.4e-07 PS=4.8e-07 $X=124520 $Y=70180 $D=1
M476 621 184 189 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.5e-14 AS=1.2e-14 PD=5e-07 PS=4.4e-07 $X=124520 $Y=71040 $D=1
M477 GND 185 621 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.2e-14 AS=1.5e-14 PD=4.4e-07 PS=5e-07 $X=124520 $Y=71440 $D=1
M478 387 182 185 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.2e-14 AS=1.2e-14 PD=4.4e-07 PS=4.4e-07 $X=124520 $Y=72300 $D=1
M479 GND 388 387 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.2e-14 AS=1.2e-14 PD=4.4e-07 PS=4.4e-07 $X=124520 $Y=73160 $D=1
M480 GND A6 388 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.2e-14 AS=1.2e-14 PD=4.4e-07 PS=4.4e-07 $X=124520 $Y=74020 $D=1
M481 GND 183 S6 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.2e-14 AS=1.2e-14 PD=4.4e-07 PS=4.4e-07 $X=124525 $Y=49225 $D=1
M482 GND 386 390 GND NMOS_VTL L=5e-08 W=1.15e-07 AD=1.61e-14 AS=1.3225e-14 PD=5.1e-07 PS=4.6e-07 $X=125060 $Y=54555 $D=1
M483 GND 386 392 GND NMOS_VTL L=5e-08 W=1.15e-07 AD=1.61e-14 AS=1.3225e-14 PD=5.1e-07 PS=4.6e-07 $X=125060 $Y=57635 $D=1
M484 GND 183 186 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.2e-14 AS=1.2e-14 PD=4.4e-07 PS=4.4e-07 $X=125385 $Y=49225 $D=1
M485 390 389 GND GND NMOS_VTL L=5e-08 W=1.15e-07 AD=1.61e-14 AS=1.61e-14 PD=5.1e-07 PS=5.1e-07 $X=125440 $Y=54555 $D=1
M486 392 389 GND GND NMOS_VTL L=5e-08 W=1.15e-07 AD=1.61e-14 AS=1.61e-14 PD=5.1e-07 PS=5.1e-07 $X=125440 $Y=57635 $D=1
M487 195 166 390 GND NMOS_VTL L=5e-08 W=1.15e-07 AD=1.61e-14 AS=1.61e-14 PD=5.1e-07 PS=5.1e-07 $X=125820 $Y=54555 $D=1
M488 196 167 392 GND NMOS_VTL L=5e-08 W=1.15e-07 AD=1.61e-14 AS=1.61e-14 PD=5.1e-07 PS=5.1e-07 $X=125820 $Y=57635 $D=1
M489 622 386 195 GND NMOS_VTL L=5e-08 W=1.15e-07 AD=1.61e-14 AS=1.61e-14 PD=5.1e-07 PS=5.1e-07 $X=126200 $Y=54555 $D=1
M490 623 386 196 GND NMOS_VTL L=5e-08 W=1.15e-07 AD=1.61e-14 AS=1.61e-14 PD=5.1e-07 PS=5.1e-07 $X=126200 $Y=57635 $D=1
M491 624 186 183 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.5e-14 AS=1.2e-14 PD=5e-07 PS=4.4e-07 $X=126245 $Y=49225 $D=1
M492 GND 389 622 GND NMOS_VTL L=5e-08 W=1.15e-07 AD=1.3225e-14 AS=1.61e-14 PD=4.6e-07 PS=5.1e-07 $X=126580 $Y=54555 $D=1
M493 GND 389 623 GND NMOS_VTL L=5e-08 W=1.15e-07 AD=1.3225e-14 AS=1.61e-14 PD=4.6e-07 PS=5.1e-07 $X=126580 $Y=57635 $D=1
M494 625 194 624 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.4e-14 AS=1.5e-14 PD=4.8e-07 PS=5e-07 $X=126645 $Y=49225 $D=1
M495 GND 192 625 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.2e-14 AS=1.4e-14 PD=4.4e-07 PS=4.8e-07 $X=127025 $Y=49225 $D=1
M496 395 386 GND GND NMOS_VTL L=5e-08 W=1e-07 AD=1.4e-14 AS=1.15e-14 PD=4.8e-07 PS=4.3e-07 $X=127300 $Y=54585 $D=1
M497 397 386 GND GND NMOS_VTL L=5e-08 W=1e-07 AD=1.4e-14 AS=1.15e-14 PD=4.8e-07 PS=4.3e-07 $X=127300 $Y=57665 $D=1
M498 GND 389 395 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.4e-14 AS=1.4e-14 PD=4.8e-07 PS=4.8e-07 $X=127680 $Y=54585 $D=1
M499 GND 389 397 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.4e-14 AS=1.4e-14 PD=4.8e-07 PS=4.8e-07 $X=127680 $Y=57665 $D=1
M500 GND RESET 194 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.2e-14 AS=1.2e-14 PD=4.4e-07 PS=4.4e-07 $X=127905 $Y=49225 $D=1
M501 395 166 GND GND NMOS_VTL L=5e-08 W=1e-07 AD=1.15e-14 AS=1.4e-14 PD=4.3e-07 PS=4.8e-07 $X=128060 $Y=54585 $D=1
M502 397 167 GND GND NMOS_VTL L=5e-08 W=1e-07 AD=1.15e-14 AS=1.4e-14 PD=4.3e-07 PS=4.8e-07 $X=128060 $Y=57665 $D=1
M503 GND 192 193 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.2e-14 AS=1.2e-14 PD=4.4e-07 PS=4.4e-07 $X=128765 $Y=49225 $D=1
M504 399 195 395 GND NMOS_VTL L=5e-08 W=9e-08 AD=1.08e-14 AS=1.125e-14 PD=4.2e-07 PS=4.3e-07 $X=128800 $Y=54585 $D=1
M505 400 196 397 GND NMOS_VTL L=5e-08 W=9e-08 AD=1.08e-14 AS=1.125e-14 PD=4.2e-07 PS=4.3e-07 $X=128800 $Y=57665 $D=1
M506 626 166 399 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.4e-14 AS=1.15e-14 PD=4.8e-07 PS=4.3e-07 $X=129530 $Y=54585 $D=1
M507 627 167 400 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.4e-14 AS=1.15e-14 PD=4.8e-07 PS=4.3e-07 $X=129530 $Y=57665 $D=1
M508 GND 18 192 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.2e-14 AS=1.2e-14 PD=4.4e-07 PS=4.4e-07 $X=129625 $Y=49225 $D=1
M509 628 386 626 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.4e-14 AS=1.4e-14 PD=4.8e-07 PS=4.8e-07 $X=129910 $Y=54585 $D=1
M510 629 386 627 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.4e-14 AS=1.4e-14 PD=4.8e-07 PS=4.8e-07 $X=129910 $Y=57665 $D=1
M511 GND 202 389 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.2e-14 AS=1.2e-14 PD=4.4e-07 PS=4.4e-07 $X=130020 $Y=62980 $D=1
M512 GND 202 201 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.2e-14 AS=1.2e-14 PD=4.4e-07 PS=4.4e-07 $X=130020 $Y=63840 $D=1
M513 630 201 202 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.5e-14 AS=1.2e-14 PD=5e-07 PS=4.4e-07 $X=130020 $Y=64700 $D=1
M514 631 199 630 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.4e-14 AS=1.5e-14 PD=4.8e-07 PS=5e-07 $X=130020 $Y=65100 $D=1
M515 GND 198 631 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.2e-14 AS=1.4e-14 PD=4.4e-07 PS=4.8e-07 $X=130020 $Y=65480 $D=1
M516 GND RESET 199 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.2e-14 AS=1.2e-14 PD=4.4e-07 PS=4.4e-07 $X=130020 $Y=66360 $D=1
M517 GND 198 197 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.2e-14 AS=1.2e-14 PD=4.4e-07 PS=4.4e-07 $X=130020 $Y=67220 $D=1
M518 GND 18 198 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.2e-14 AS=1.2e-14 PD=4.4e-07 PS=4.4e-07 $X=130020 $Y=68080 $D=1
M519 203 197 202 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.2e-14 AS=1.2e-14 PD=4.4e-07 PS=4.4e-07 $X=130020 $Y=68940 $D=1
M520 632 197 GND GND NMOS_VTL L=5e-08 W=1e-07 AD=1.4e-14 AS=1.2e-14 PD=4.8e-07 PS=4.4e-07 $X=130020 $Y=69800 $D=1
M521 200 203 632 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.2e-14 AS=1.4e-14 PD=4.4e-07 PS=4.8e-07 $X=130020 $Y=70180 $D=1
M522 633 199 203 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.5e-14 AS=1.2e-14 PD=5e-07 PS=4.4e-07 $X=130020 $Y=71040 $D=1
M523 GND 200 633 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.2e-14 AS=1.5e-14 PD=4.4e-07 PS=5e-07 $X=130020 $Y=71440 $D=1
M524 401 198 200 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.2e-14 AS=1.2e-14 PD=4.4e-07 PS=4.4e-07 $X=130020 $Y=72300 $D=1
M525 GND 402 401 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.2e-14 AS=1.2e-14 PD=4.4e-07 PS=4.4e-07 $X=130020 $Y=73160 $D=1
M526 GND B6 402 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.2e-14 AS=1.2e-14 PD=4.4e-07 PS=4.4e-07 $X=130020 $Y=74020 $D=1
M527 GND 389 628 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.15e-14 AS=1.4e-14 PD=4.3e-07 PS=4.8e-07 $X=130290 $Y=54585 $D=1
M528 GND 389 629 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.15e-14 AS=1.4e-14 PD=4.3e-07 PS=4.8e-07 $X=130290 $Y=57665 $D=1
M529 204 193 183 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.2e-14 AS=1.2e-14 PD=4.4e-07 PS=4.4e-07 $X=130485 $Y=49225 $D=1
M530 634 193 GND GND NMOS_VTL L=5e-08 W=1e-07 AD=1.4e-14 AS=1.2e-14 PD=4.8e-07 PS=4.4e-07 $X=131345 $Y=49225 $D=1
M531 210 399 GND GND NMOS_VTL L=5e-08 W=1e-07 AD=1.2e-14 AS=1.2e-14 PD=4.4e-07 PS=4.4e-07 $X=131395 $Y=55135 $D=1
M532 404 121 GND GND NMOS_VTL L=5e-08 W=1e-07 AD=1.35e-14 AS=1.15e-14 PD=4.7e-07 PS=4.3e-07 $X=131420 $Y=57305 $D=1
M533 207 204 634 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.2e-14 AS=1.4e-14 PD=4.4e-07 PS=4.8e-07 $X=131725 $Y=49225 $D=1
M534 209 404 208 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.4e-14 AS=1.2e-14 PD=4.8e-07 PS=4.4e-07 $X=132190 $Y=57305 $D=1
M535 GND 400 208 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.2e-14 AS=1.2e-14 PD=4.4e-07 PS=4.4e-07 $X=132400 $Y=58455 $D=1
M536 210 121 209 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.15e-14 AS=1.4e-14 PD=4.3e-07 PS=4.8e-07 $X=132570 $Y=57305 $D=1
M537 635 194 204 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.5e-14 AS=1.2e-14 PD=5e-07 PS=4.4e-07 $X=132585 $Y=49225 $D=1
M538 GND 207 635 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.2e-14 AS=1.5e-14 PD=4.4e-07 PS=5e-07 $X=132985 $Y=49225 $D=1
M539 405 192 207 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.2e-14 AS=1.2e-14 PD=4.4e-07 PS=4.4e-07 $X=133845 $Y=49225 $D=1
M540 GND 406 405 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.2e-14 AS=1.2e-14 PD=4.4e-07 PS=4.4e-07 $X=134705 $Y=49225 $D=1
M541 GND 209 406 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.2e-14 AS=1.2e-14 PD=4.4e-07 PS=4.4e-07 $X=135565 $Y=49225 $D=1
M542 GND 410 409 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.2e-14 AS=1.2e-14 PD=4.4e-07 PS=4.4e-07 $X=136225 $Y=61795 $D=1
M543 GND 216 410 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.2e-14 AS=1.2e-14 PD=4.4e-07 PS=4.4e-07 $X=136225 $Y=62980 $D=1
M544 GND 216 215 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.2e-14 AS=1.2e-14 PD=4.4e-07 PS=4.4e-07 $X=136225 $Y=63840 $D=1
M545 636 215 216 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.5e-14 AS=1.2e-14 PD=5e-07 PS=4.4e-07 $X=136225 $Y=64700 $D=1
M546 637 213 636 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.4e-14 AS=1.5e-14 PD=4.8e-07 PS=5e-07 $X=136225 $Y=65100 $D=1
M547 GND 212 637 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.2e-14 AS=1.4e-14 PD=4.4e-07 PS=4.8e-07 $X=136225 $Y=65480 $D=1
M548 GND RESET 213 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.2e-14 AS=1.2e-14 PD=4.4e-07 PS=4.4e-07 $X=136225 $Y=66360 $D=1
M549 GND 212 211 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.2e-14 AS=1.2e-14 PD=4.4e-07 PS=4.4e-07 $X=136225 $Y=67220 $D=1
M550 GND 18 212 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.2e-14 AS=1.2e-14 PD=4.4e-07 PS=4.4e-07 $X=136225 $Y=68080 $D=1
M551 217 211 216 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.2e-14 AS=1.2e-14 PD=4.4e-07 PS=4.4e-07 $X=136225 $Y=68940 $D=1
M552 638 211 GND GND NMOS_VTL L=5e-08 W=1e-07 AD=1.4e-14 AS=1.2e-14 PD=4.8e-07 PS=4.4e-07 $X=136225 $Y=69800 $D=1
M553 214 217 638 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.2e-14 AS=1.4e-14 PD=4.4e-07 PS=4.8e-07 $X=136225 $Y=70180 $D=1
M554 639 213 217 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.5e-14 AS=1.2e-14 PD=5e-07 PS=4.4e-07 $X=136225 $Y=71040 $D=1
M555 GND 214 639 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.2e-14 AS=1.5e-14 PD=4.4e-07 PS=5e-07 $X=136225 $Y=71440 $D=1
M556 411 212 214 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.2e-14 AS=1.2e-14 PD=4.4e-07 PS=4.4e-07 $X=136225 $Y=72300 $D=1
M557 GND 412 411 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.2e-14 AS=1.2e-14 PD=4.4e-07 PS=4.4e-07 $X=136225 $Y=73160 $D=1
M558 GND A7 412 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.2e-14 AS=1.2e-14 PD=4.4e-07 PS=4.4e-07 $X=136225 $Y=74020 $D=1
M559 GND 409 414 GND NMOS_VTL L=5e-08 W=1.15e-07 AD=1.61e-14 AS=1.3225e-14 PD=5.1e-07 PS=4.6e-07 $X=136860 $Y=54555 $D=1
M560 GND 409 416 GND NMOS_VTL L=5e-08 W=1.15e-07 AD=1.61e-14 AS=1.3225e-14 PD=5.1e-07 PS=4.6e-07 $X=136860 $Y=57635 $D=1
M561 GND 218 S7 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.2e-14 AS=1.2e-14 PD=4.4e-07 PS=4.4e-07 $X=136905 $Y=49225 $D=1
M562 414 413 GND GND NMOS_VTL L=5e-08 W=1.15e-07 AD=1.61e-14 AS=1.61e-14 PD=5.1e-07 PS=5.1e-07 $X=137240 $Y=54555 $D=1
M563 416 413 GND GND NMOS_VTL L=5e-08 W=1.15e-07 AD=1.61e-14 AS=1.61e-14 PD=5.1e-07 PS=5.1e-07 $X=137240 $Y=57635 $D=1
M564 225 195 414 GND NMOS_VTL L=5e-08 W=1.15e-07 AD=1.61e-14 AS=1.61e-14 PD=5.1e-07 PS=5.1e-07 $X=137620 $Y=54555 $D=1
M565 226 196 416 GND NMOS_VTL L=5e-08 W=1.15e-07 AD=1.61e-14 AS=1.61e-14 PD=5.1e-07 PS=5.1e-07 $X=137620 $Y=57635 $D=1
M566 GND 218 220 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.2e-14 AS=1.2e-14 PD=4.4e-07 PS=4.4e-07 $X=137765 $Y=49225 $D=1
M567 640 409 225 GND NMOS_VTL L=5e-08 W=1.15e-07 AD=1.61e-14 AS=1.61e-14 PD=5.1e-07 PS=5.1e-07 $X=138000 $Y=54555 $D=1
M568 641 409 226 GND NMOS_VTL L=5e-08 W=1.15e-07 AD=1.61e-14 AS=1.61e-14 PD=5.1e-07 PS=5.1e-07 $X=138000 $Y=57635 $D=1
M569 GND 413 640 GND NMOS_VTL L=5e-08 W=1.15e-07 AD=1.3225e-14 AS=1.61e-14 PD=4.6e-07 PS=5.1e-07 $X=138380 $Y=54555 $D=1
M570 GND 413 641 GND NMOS_VTL L=5e-08 W=1.15e-07 AD=1.3225e-14 AS=1.61e-14 PD=4.6e-07 PS=5.1e-07 $X=138380 $Y=57635 $D=1
M571 642 220 218 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.5e-14 AS=1.2e-14 PD=5e-07 PS=4.4e-07 $X=138625 $Y=49225 $D=1
M572 643 224 642 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.4e-14 AS=1.5e-14 PD=4.8e-07 PS=5e-07 $X=139025 $Y=49225 $D=1
M573 419 409 GND GND NMOS_VTL L=5e-08 W=1e-07 AD=1.4e-14 AS=1.15e-14 PD=4.8e-07 PS=4.3e-07 $X=139100 $Y=54585 $D=1
M574 421 409 GND GND NMOS_VTL L=5e-08 W=1e-07 AD=1.4e-14 AS=1.15e-14 PD=4.8e-07 PS=4.3e-07 $X=139100 $Y=57665 $D=1
M575 GND 222 643 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.2e-14 AS=1.4e-14 PD=4.4e-07 PS=4.8e-07 $X=139405 $Y=49225 $D=1
M576 GND 413 419 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.4e-14 AS=1.4e-14 PD=4.8e-07 PS=4.8e-07 $X=139480 $Y=54585 $D=1
M577 GND 413 421 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.4e-14 AS=1.4e-14 PD=4.8e-07 PS=4.8e-07 $X=139480 $Y=57665 $D=1
M578 419 195 GND GND NMOS_VTL L=5e-08 W=1e-07 AD=1.15e-14 AS=1.4e-14 PD=4.3e-07 PS=4.8e-07 $X=139860 $Y=54585 $D=1
M579 421 196 GND GND NMOS_VTL L=5e-08 W=1e-07 AD=1.15e-14 AS=1.4e-14 PD=4.3e-07 PS=4.8e-07 $X=139860 $Y=57665 $D=1
M580 GND RESET 224 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.2e-14 AS=1.2e-14 PD=4.4e-07 PS=4.4e-07 $X=140285 $Y=49225 $D=1
M581 423 225 419 GND NMOS_VTL L=5e-08 W=9e-08 AD=1.08e-14 AS=1.125e-14 PD=4.2e-07 PS=4.3e-07 $X=140600 $Y=54585 $D=1
M582 236 226 421 GND NMOS_VTL L=5e-08 W=9e-08 AD=1.08e-14 AS=1.125e-14 PD=4.2e-07 PS=4.3e-07 $X=140600 $Y=57665 $D=1
M583 GND 222 223 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.2e-14 AS=1.2e-14 PD=4.4e-07 PS=4.4e-07 $X=141145 $Y=49225 $D=1
M584 644 195 423 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.4e-14 AS=1.15e-14 PD=4.8e-07 PS=4.3e-07 $X=141330 $Y=54585 $D=1
M585 645 196 236 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.4e-14 AS=1.15e-14 PD=4.8e-07 PS=4.3e-07 $X=141330 $Y=57665 $D=1
M586 650 409 644 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.4e-14 AS=1.4e-14 PD=4.8e-07 PS=4.8e-07 $X=141710 $Y=54585 $D=1
M587 651 409 645 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.4e-14 AS=1.4e-14 PD=4.8e-07 PS=4.8e-07 $X=141710 $Y=57665 $D=1
M588 GND 424 413 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.2e-14 AS=1.2e-14 PD=4.4e-07 PS=4.4e-07 $X=141745 $Y=61795 $D=1
M589 GND 232 424 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.2e-14 AS=1.2e-14 PD=4.4e-07 PS=4.4e-07 $X=141745 $Y=62980 $D=1
M590 GND 232 231 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.2e-14 AS=1.2e-14 PD=4.4e-07 PS=4.4e-07 $X=141745 $Y=63840 $D=1
M591 646 231 232 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.5e-14 AS=1.2e-14 PD=5e-07 PS=4.4e-07 $X=141745 $Y=64700 $D=1
M592 647 229 646 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.4e-14 AS=1.5e-14 PD=4.8e-07 PS=5e-07 $X=141745 $Y=65100 $D=1
M593 GND 228 647 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.2e-14 AS=1.4e-14 PD=4.4e-07 PS=4.8e-07 $X=141745 $Y=65480 $D=1
M594 GND RESET 229 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.2e-14 AS=1.2e-14 PD=4.4e-07 PS=4.4e-07 $X=141745 $Y=66360 $D=1
M595 GND 228 227 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.2e-14 AS=1.2e-14 PD=4.4e-07 PS=4.4e-07 $X=141745 $Y=67220 $D=1
M596 GND 18 228 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.2e-14 AS=1.2e-14 PD=4.4e-07 PS=4.4e-07 $X=141745 $Y=68080 $D=1
M597 233 227 232 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.2e-14 AS=1.2e-14 PD=4.4e-07 PS=4.4e-07 $X=141745 $Y=68940 $D=1
M598 648 227 GND GND NMOS_VTL L=5e-08 W=1e-07 AD=1.4e-14 AS=1.2e-14 PD=4.8e-07 PS=4.4e-07 $X=141745 $Y=69800 $D=1
M599 230 233 648 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.2e-14 AS=1.4e-14 PD=4.4e-07 PS=4.8e-07 $X=141745 $Y=70180 $D=1
M600 649 229 233 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.5e-14 AS=1.2e-14 PD=5e-07 PS=4.4e-07 $X=141745 $Y=71040 $D=1
M601 GND 230 649 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.2e-14 AS=1.5e-14 PD=4.4e-07 PS=5e-07 $X=141745 $Y=71440 $D=1
M602 425 228 230 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.2e-14 AS=1.2e-14 PD=4.4e-07 PS=4.4e-07 $X=141745 $Y=72300 $D=1
M603 GND 426 425 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.2e-14 AS=1.2e-14 PD=4.4e-07 PS=4.4e-07 $X=141745 $Y=73160 $D=1
M604 GND B7 426 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.2e-14 AS=1.2e-14 PD=4.4e-07 PS=4.4e-07 $X=141745 $Y=74020 $D=1
M605 GND 18 222 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.2e-14 AS=1.2e-14 PD=4.4e-07 PS=4.4e-07 $X=142005 $Y=49225 $D=1
M606 GND 413 650 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.15e-14 AS=1.4e-14 PD=4.3e-07 PS=4.8e-07 $X=142090 $Y=54585 $D=1
M607 GND 413 651 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.15e-14 AS=1.4e-14 PD=4.3e-07 PS=4.8e-07 $X=142090 $Y=57665 $D=1
M608 235 223 218 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.2e-14 AS=1.2e-14 PD=4.4e-07 PS=4.4e-07 $X=142865 $Y=49225 $D=1
M609 429 121 GND GND NMOS_VTL L=5e-08 W=1e-07 AD=1.35e-14 AS=1.15e-14 PD=4.7e-07 PS=4.3e-07 $X=143220 $Y=57305 $D=1
M610 652 223 GND GND NMOS_VTL L=5e-08 W=1e-07 AD=1.4e-14 AS=1.2e-14 PD=4.8e-07 PS=4.4e-07 $X=143725 $Y=49225 $D=1
M611 237 429 236 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.4e-14 AS=1.2e-14 PD=4.8e-07 PS=4.4e-07 $X=143990 $Y=57305 $D=1
M612 238 235 652 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.2e-14 AS=1.4e-14 PD=4.4e-07 PS=4.8e-07 $X=144105 $Y=49225 $D=1
M613 239 121 237 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.15e-14 AS=1.4e-14 PD=4.3e-07 PS=4.8e-07 $X=144370 $Y=57305 $D=1
M614 653 224 235 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.5e-14 AS=1.2e-14 PD=5e-07 PS=4.4e-07 $X=144965 $Y=49225 $D=1
M615 GND 238 653 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.2e-14 AS=1.5e-14 PD=4.4e-07 PS=5e-07 $X=145365 $Y=49225 $D=1
M616 431 222 238 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.2e-14 AS=1.2e-14 PD=4.4e-07 PS=4.4e-07 $X=146225 $Y=49225 $D=1
M617 430 121 GND GND NMOS_VTL L=5e-08 W=1e-07 AD=1.35e-14 AS=1.15e-14 PD=4.7e-07 PS=4.3e-07 $X=146325 $Y=57280 $D=1
M618 GND 432 431 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.2e-14 AS=1.2e-14 PD=4.4e-07 PS=4.4e-07 $X=147085 $Y=49225 $D=1
M619 VDD 430 226 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.4e-14 AS=1.2e-14 PD=4.8e-07 PS=4.4e-07 $X=147095 $Y=57280 $D=1
M620 225 121 VDD GND NMOS_VTL L=5e-08 W=1e-07 AD=1.15e-14 AS=1.4e-14 PD=4.3e-07 PS=4.8e-07 $X=147475 $Y=57280 $D=1
M621 GND 237 432 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.2e-14 AS=1.2e-14 PD=4.4e-07 PS=4.4e-07 $X=147945 $Y=49225 $D=1
M622 435 VDD GND GND NMOS_VTL L=5e-08 W=1e-07 AD=1.2e-14 AS=1.2e-14 PD=4.4e-07 PS=4.4e-07 $X=150115 $Y=57685 $D=1
M623 436 435 GND GND NMOS_VTL L=5e-08 W=1e-07 AD=1.2e-14 AS=1.2e-14 PD=4.4e-07 PS=4.4e-07 $X=150115 $Y=58545 $D=1
M624 246 244 436 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.2e-14 AS=1.2e-14 PD=4.4e-07 PS=4.4e-07 $X=150115 $Y=59405 $D=1
M625 654 246 GND GND NMOS_VTL L=5e-08 W=1e-07 AD=1.5e-14 AS=1.2e-14 PD=5e-07 PS=4.4e-07 $X=150115 $Y=60265 $D=1
M626 247 243 654 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.2e-14 AS=1.5e-14 PD=4.4e-07 PS=5e-07 $X=150115 $Y=60665 $D=1
M627 655 247 246 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.4e-14 AS=1.2e-14 PD=4.8e-07 PS=4.4e-07 $X=150115 $Y=61525 $D=1
M628 GND 240 655 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.2e-14 AS=1.4e-14 PD=4.4e-07 PS=4.8e-07 $X=150115 $Y=61905 $D=1
M629 242 240 247 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.2e-14 AS=1.2e-14 PD=4.4e-07 PS=4.4e-07 $X=150115 $Y=62765 $D=1
M630 244 18 GND GND NMOS_VTL L=5e-08 W=1e-07 AD=1.2e-14 AS=1.2e-14 PD=4.4e-07 PS=4.4e-07 $X=150115 $Y=63625 $D=1
M631 240 244 GND GND NMOS_VTL L=5e-08 W=1e-07 AD=1.2e-14 AS=1.2e-14 PD=4.4e-07 PS=4.4e-07 $X=150115 $Y=64485 $D=1
M632 243 RESET GND GND NMOS_VTL L=5e-08 W=1e-07 AD=1.2e-14 AS=1.2e-14 PD=4.4e-07 PS=4.4e-07 $X=150115 $Y=65345 $D=1
M633 656 244 GND GND NMOS_VTL L=5e-08 W=1e-07 AD=1.4e-14 AS=1.2e-14 PD=4.8e-07 PS=4.4e-07 $X=150115 $Y=66225 $D=1
M634 657 243 656 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.5e-14 AS=1.4e-14 PD=5e-07 PS=4.8e-07 $X=150115 $Y=66605 $D=1
M635 242 241 657 GND NMOS_VTL L=5e-08 W=1e-07 AD=1.2e-14 AS=1.5e-14 PD=4.4e-07 PS=5e-07 $X=150115 $Y=67005 $D=1
M636 241 242 GND GND NMOS_VTL L=5e-08 W=1e-07 AD=1.2e-14 AS=1.2e-14 PD=4.4e-07 PS=4.4e-07 $X=150115 $Y=67865 $D=1
M637 434 242 GND GND NMOS_VTL L=5e-08 W=1e-07 AD=1.2e-14 AS=1.2e-14 PD=4.4e-07 PS=4.4e-07 $X=150115 $Y=68725 $D=1
M638 270 5 S0 270 PMOS_VTL L=5e-08 W=1.6e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 $X=49850 $Y=50125 $D=0
M639 270 5 6 270 PMOS_VTL L=5e-08 W=1.6e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 $X=50710 $Y=50125 $D=0
M640 VDD 249 254 VDD PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=2.07e-14 PD=6.4e-07 PS=5.9e-07 $X=50990 $Y=55935 $D=0
M641 VDD 249 256 VDD PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=2.07e-14 PD=6.4e-07 PS=5.9e-07 $X=50990 $Y=58855 $D=0
M642 VDD 10 249 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 $X=51350 $Y=62980 $D=0
M643 VDD 10 9 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 $X=51350 $Y=63840 $D=0
M644 10 9 13 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=2.4e-14 AS=1.92e-14 PD=6.2e-07 PS=5.6e-07 $X=51350 $Y=64700 $D=0
M645 13 7 10 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=2.4e-14 AS=2.4e-14 PD=6.2e-07 PS=6.2e-07 $X=51350 $Y=65100 $D=0
M646 VDD 3 13 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=1.92e-14 AS=2.4e-14 PD=5.6e-07 PS=6.2e-07 $X=51350 $Y=65500 $D=0
M647 VDD RESET 7 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 $X=51350 $Y=66360 $D=0
M648 VDD 4 3 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 $X=51350 $Y=67220 $D=0
M649 VDD 18 4 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 $X=51350 $Y=68080 $D=0
M650 11 4 10 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 $X=51350 $Y=68940 $D=0
M651 437 4 VDD VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=2.24e-14 AS=1.92e-14 PD=6e-07 PS=5.6e-07 $X=51350 $Y=69800 $D=0
M652 8 11 437 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=1.92e-14 AS=2.24e-14 PD=5.6e-07 PS=6e-07 $X=51350 $Y=70180 $D=0
M653 11 7 VDD VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=2.4e-14 AS=1.92e-14 PD=6.2e-07 PS=5.6e-07 $X=51350 $Y=71040 $D=0
M654 VDD 8 11 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=1.92e-14 AS=2.4e-14 PD=5.6e-07 PS=6.2e-07 $X=51350 $Y=71440 $D=0
M655 250 3 8 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 $X=51350 $Y=72300 $D=0
M656 VDD 251 250 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 $X=51350 $Y=73160 $D=0
M657 VDD A0 251 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 $X=51350 $Y=74020 $D=0
M658 254 252 VDD VDD PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=2.52e-14 PD=6.4e-07 PS=6.4e-07 $X=51370 $Y=55935 $D=0
M659 256 252 VDD VDD PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=2.52e-14 PD=6.4e-07 PS=6.4e-07 $X=51370 $Y=58855 $D=0
M660 5 6 12 270 PMOS_VTL L=5e-08 W=1.6e-07 AD=2.4e-14 AS=1.92e-14 PD=6.2e-07 PS=5.6e-07 $X=51570 $Y=50125 $D=0
M661 19 VDD 254 VDD PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=2.52e-14 PD=6.4e-07 PS=6.4e-07 $X=51750 $Y=55935 $D=0
M662 20 GND 256 VDD PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=2.52e-14 PD=6.4e-07 PS=6.4e-07 $X=51750 $Y=58855 $D=0
M663 12 17 5 270 PMOS_VTL L=5e-08 W=1.6e-07 AD=2.4e-14 AS=2.4e-14 PD=6.2e-07 PS=6.2e-07 $X=51970 $Y=50125 $D=0
M664 438 249 19 VDD PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=2.52e-14 PD=6.4e-07 PS=6.4e-07 $X=52130 $Y=55935 $D=0
M665 439 249 20 VDD PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=2.52e-14 PD=6.4e-07 PS=6.4e-07 $X=52130 $Y=58855 $D=0
M666 270 15 12 270 PMOS_VTL L=5e-08 W=1.6e-07 AD=1.92e-14 AS=2.4e-14 PD=5.6e-07 PS=6.2e-07 $X=52370 $Y=50125 $D=0
M667 VDD 252 438 VDD PMOS_VTL L=5e-08 W=1.8e-07 AD=2.07e-14 AS=2.52e-14 PD=5.9e-07 PS=6.4e-07 $X=52510 $Y=55935 $D=0
M668 VDD 252 439 VDD PMOS_VTL L=5e-08 W=1.8e-07 AD=2.07e-14 AS=2.52e-14 PD=5.9e-07 PS=6.4e-07 $X=52510 $Y=58855 $D=0
M669 270 RESET 17 270 PMOS_VTL L=5e-08 W=1.6e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 $X=53230 $Y=50125 $D=0
M670 259 249 VDD VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=2.24e-14 AS=1.84e-14 PD=6e-07 PS=5.5e-07 $X=53230 $Y=55935 $D=0
M671 261 249 VDD VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=2.24e-14 AS=1.84e-14 PD=6e-07 PS=5.5e-07 $X=53230 $Y=58855 $D=0
M672 VDD 252 259 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=2.24e-14 AS=2.24e-14 PD=6e-07 PS=6e-07 $X=53610 $Y=55935 $D=0
M673 VDD 252 261 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=2.24e-14 AS=2.24e-14 PD=6e-07 PS=6e-07 $X=53610 $Y=58855 $D=0
M674 259 VDD VDD VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=1.84e-14 AS=2.24e-14 PD=5.5e-07 PS=6e-07 $X=53990 $Y=55935 $D=0
M675 261 GND VDD VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=1.84e-14 AS=2.24e-14 PD=5.5e-07 PS=6e-07 $X=53990 $Y=58855 $D=0
M676 270 14 15 270 PMOS_VTL L=5e-08 W=1.6e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 $X=54090 $Y=50125 $D=0
M677 262 19 259 VDD PMOS_VTL L=5e-08 W=1.4e-07 AD=1.68e-14 AS=1.75e-14 PD=5.2e-07 PS=5.3e-07 $X=54730 $Y=55935 $D=0
M678 263 20 261 VDD PMOS_VTL L=5e-08 W=1.4e-07 AD=1.68e-14 AS=1.75e-14 PD=5.2e-07 PS=5.3e-07 $X=54730 $Y=58855 $D=0
M679 270 18 14 270 PMOS_VTL L=5e-08 W=1.6e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 $X=54950 $Y=50125 $D=0
M680 440 VDD 262 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=2.24e-14 AS=1.84e-14 PD=6e-07 PS=5.5e-07 $X=55460 $Y=55935 $D=0
M681 441 GND 263 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=2.24e-14 AS=1.84e-14 PD=6e-07 PS=5.5e-07 $X=55460 $Y=58855 $D=0
M682 23 14 5 270 PMOS_VTL L=5e-08 W=1.6e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 $X=55810 $Y=50125 $D=0
M683 442 249 440 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=2.24e-14 AS=2.24e-14 PD=6e-07 PS=6e-07 $X=55840 $Y=55935 $D=0
M684 443 249 441 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=2.24e-14 AS=2.24e-14 PD=6e-07 PS=6e-07 $X=55840 $Y=58855 $D=0
M685 VDD 252 442 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=1.84e-14 AS=2.24e-14 PD=5.5e-07 PS=6e-07 $X=56220 $Y=55935 $D=0
M686 VDD 252 443 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=1.84e-14 AS=2.24e-14 PD=5.5e-07 PS=6e-07 $X=56220 $Y=58855 $D=0
M687 444 14 270 270 PMOS_VTL L=5e-08 W=1.6e-07 AD=2.24e-14 AS=1.92e-14 PD=6e-07 PS=5.6e-07 $X=56670 $Y=50125 $D=0
M688 VDD 27 252 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 $X=56850 $Y=62980 $D=0
M689 VDD 27 26 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 $X=56850 $Y=63840 $D=0
M690 27 26 29 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=2.4e-14 AS=1.92e-14 PD=6.2e-07 PS=5.6e-07 $X=56850 $Y=64700 $D=0
M691 29 24 27 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=2.4e-14 AS=2.4e-14 PD=6.2e-07 PS=6.2e-07 $X=56850 $Y=65100 $D=0
M692 VDD 21 29 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=1.92e-14 AS=2.4e-14 PD=5.6e-07 PS=6.2e-07 $X=56850 $Y=65500 $D=0
M693 VDD RESET 24 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 $X=56850 $Y=66360 $D=0
M694 VDD 22 21 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 $X=56850 $Y=67220 $D=0
M695 VDD 18 22 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 $X=56850 $Y=68080 $D=0
M696 28 22 27 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 $X=56850 $Y=68940 $D=0
M697 445 22 VDD VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=2.24e-14 AS=1.92e-14 PD=6e-07 PS=5.6e-07 $X=56850 $Y=69800 $D=0
M698 25 28 445 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=1.92e-14 AS=2.24e-14 PD=5.6e-07 PS=6e-07 $X=56850 $Y=70180 $D=0
M699 28 24 VDD VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=2.4e-14 AS=1.92e-14 PD=6.2e-07 PS=5.6e-07 $X=56850 $Y=71040 $D=0
M700 VDD 25 28 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=1.92e-14 AS=2.4e-14 PD=5.6e-07 PS=6.2e-07 $X=56850 $Y=71440 $D=0
M701 264 21 25 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 $X=56850 $Y=72300 $D=0
M702 VDD 265 264 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 $X=56850 $Y=73160 $D=0
M703 VDD B0 265 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 $X=56850 $Y=74020 $D=0
M704 30 23 444 270 PMOS_VTL L=5e-08 W=1.6e-07 AD=1.92e-14 AS=2.24e-14 PD=5.6e-07 PS=6e-07 $X=57050 $Y=50125 $D=0
M705 VDD 263 31 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 $X=57320 $Y=58455 $D=0
M706 267 GND VDD VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=1.84e-14 AS=1.84e-14 PD=5.5e-07 PS=5.5e-07 $X=57350 $Y=56315 $D=0
M707 23 17 270 270 PMOS_VTL L=5e-08 W=1.6e-07 AD=2.4e-14 AS=1.92e-14 PD=6.2e-07 PS=5.6e-07 $X=57910 $Y=50125 $D=0
M708 32 GND 31 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=2.24e-14 AS=1.84e-14 PD=6e-07 PS=5.5e-07 $X=58120 $Y=56315 $D=0
M709 33 262 VDD VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 $X=58215 $Y=55295 $D=0
M710 270 30 23 270 PMOS_VTL L=5e-08 W=1.6e-07 AD=1.92e-14 AS=2.4e-14 PD=5.6e-07 PS=6.2e-07 $X=58310 $Y=50125 $D=0
M711 33 267 32 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=1.84e-14 AS=2.24e-14 PD=5.5e-07 PS=6e-07 $X=58500 $Y=56315 $D=0
M712 268 15 30 270 PMOS_VTL L=5e-08 W=1.6e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 $X=59170 $Y=50125 $D=0
M713 270 269 268 270 PMOS_VTL L=5e-08 W=1.6e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 $X=60030 $Y=50125 $D=0
M714 270 32 269 270 PMOS_VTL L=5e-08 W=1.6e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 $X=60890 $Y=50125 $D=0
M715 291 36 S1 291 PMOS_VTL L=5e-08 W=1.6e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 $X=62115 $Y=50125 $D=0
M716 VDD VDD 277 VDD PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=2.07e-14 PD=6.4e-07 PS=5.9e-07 $X=62790 $Y=55935 $D=0
M717 VDD VDD VDD VDD PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=2.07e-14 PD=6.4e-07 PS=5.9e-07 $X=62790 $Y=59015 $D=0
M718 291 36 39 291 PMOS_VTL L=5e-08 W=1.6e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 $X=62975 $Y=50125 $D=0
M719 VDD 272 VDD VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 $X=63045 $Y=61790 $D=0
M720 VDD 41 272 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 $X=63055 $Y=62975 $D=0
M721 VDD 41 40 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 $X=63055 $Y=63835 $D=0
M722 41 40 43 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=2.4e-14 AS=1.92e-14 PD=6.2e-07 PS=5.6e-07 $X=63055 $Y=64695 $D=0
M723 43 37 41 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=2.4e-14 AS=2.4e-14 PD=6.2e-07 PS=6.2e-07 $X=63055 $Y=65095 $D=0
M724 VDD 34 43 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=1.92e-14 AS=2.4e-14 PD=5.6e-07 PS=6.2e-07 $X=63055 $Y=65495 $D=0
M725 VDD RESET 37 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 $X=63055 $Y=66355 $D=0
M726 VDD 35 34 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 $X=63055 $Y=67215 $D=0
M727 VDD 18 35 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 $X=63055 $Y=68075 $D=0
M728 42 35 41 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 $X=63055 $Y=68935 $D=0
M729 446 35 VDD VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=2.24e-14 AS=1.92e-14 PD=6e-07 PS=5.6e-07 $X=63055 $Y=69795 $D=0
M730 38 42 446 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=1.92e-14 AS=2.24e-14 PD=5.6e-07 PS=6e-07 $X=63055 $Y=70175 $D=0
M731 42 37 VDD VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=2.4e-14 AS=1.92e-14 PD=6.2e-07 PS=5.6e-07 $X=63055 $Y=71035 $D=0
M732 VDD 38 42 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=1.92e-14 AS=2.4e-14 PD=5.6e-07 PS=6.2e-07 $X=63055 $Y=71435 $D=0
M733 273 34 38 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 $X=63055 $Y=72295 $D=0
M734 VDD 274 273 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 $X=63055 $Y=73155 $D=0
M735 VDD A1 274 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 $X=63055 $Y=74015 $D=0
M736 277 275 VDD VDD PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=2.52e-14 PD=6.4e-07 PS=6.4e-07 $X=63170 $Y=55935 $D=0
M737 VDD 275 VDD VDD PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=2.52e-14 PD=6.4e-07 PS=6.4e-07 $X=63170 $Y=59015 $D=0
M738 48 19 277 VDD PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=2.52e-14 PD=6.4e-07 PS=6.4e-07 $X=63550 $Y=55935 $D=0
M739 49 20 VDD VDD PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=2.52e-14 PD=6.4e-07 PS=6.4e-07 $X=63550 $Y=59015 $D=0
M740 36 39 44 291 PMOS_VTL L=5e-08 W=1.6e-07 AD=2.4e-14 AS=1.92e-14 PD=6.2e-07 PS=5.6e-07 $X=63835 $Y=50125 $D=0
M741 447 VDD 48 VDD PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=2.52e-14 PD=6.4e-07 PS=6.4e-07 $X=63930 $Y=55935 $D=0
M742 448 VDD 49 VDD PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=2.52e-14 PD=6.4e-07 PS=6.4e-07 $X=63930 $Y=59015 $D=0
M743 44 47 36 291 PMOS_VTL L=5e-08 W=1.6e-07 AD=2.4e-14 AS=2.4e-14 PD=6.2e-07 PS=6.2e-07 $X=64235 $Y=50125 $D=0
M744 VDD 275 447 VDD PMOS_VTL L=5e-08 W=1.8e-07 AD=2.07e-14 AS=2.52e-14 PD=5.9e-07 PS=6.4e-07 $X=64310 $Y=55935 $D=0
M745 VDD 275 448 VDD PMOS_VTL L=5e-08 W=1.8e-07 AD=2.07e-14 AS=2.52e-14 PD=5.9e-07 PS=6.4e-07 $X=64310 $Y=59015 $D=0
M746 291 46 44 291 PMOS_VTL L=5e-08 W=1.6e-07 AD=1.92e-14 AS=2.4e-14 PD=5.6e-07 PS=6.2e-07 $X=64635 $Y=50125 $D=0
M747 281 VDD VDD VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=2.24e-14 AS=1.84e-14 PD=6e-07 PS=5.5e-07 $X=65030 $Y=55935 $D=0
M748 283 VDD VDD VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=2.24e-14 AS=1.84e-14 PD=6e-07 PS=5.5e-07 $X=65030 $Y=59015 $D=0
M749 VDD 275 281 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=2.24e-14 AS=2.24e-14 PD=6e-07 PS=6e-07 $X=65410 $Y=55935 $D=0
M750 VDD 275 283 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=2.24e-14 AS=2.24e-14 PD=6e-07 PS=6e-07 $X=65410 $Y=59015 $D=0
M751 291 RESET 47 291 PMOS_VTL L=5e-08 W=1.6e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 $X=65495 $Y=50125 $D=0
M752 281 19 VDD VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=1.84e-14 AS=2.24e-14 PD=5.5e-07 PS=6e-07 $X=65790 $Y=55935 $D=0
M753 283 20 VDD VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=1.84e-14 AS=2.24e-14 PD=5.5e-07 PS=6e-07 $X=65790 $Y=59015 $D=0
M754 291 45 46 291 PMOS_VTL L=5e-08 W=1.6e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 $X=66355 $Y=50125 $D=0
M755 62 48 281 VDD PMOS_VTL L=5e-08 W=1.4e-07 AD=1.68e-14 AS=1.75e-14 PD=5.2e-07 PS=5.3e-07 $X=66530 $Y=55935 $D=0
M756 60 49 283 VDD PMOS_VTL L=5e-08 W=1.4e-07 AD=1.68e-14 AS=1.75e-14 PD=5.2e-07 PS=5.3e-07 $X=66530 $Y=59015 $D=0
M757 291 18 45 291 PMOS_VTL L=5e-08 W=1.6e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 $X=67215 $Y=50125 $D=0
M758 449 19 62 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=2.24e-14 AS=1.84e-14 PD=6e-07 PS=5.5e-07 $X=67260 $Y=55935 $D=0
M759 450 20 60 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=2.24e-14 AS=1.84e-14 PD=6e-07 PS=5.5e-07 $X=67260 $Y=59015 $D=0
M760 451 VDD 449 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=2.24e-14 AS=2.24e-14 PD=6e-07 PS=6e-07 $X=67640 $Y=55935 $D=0
M761 452 VDD 450 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=2.24e-14 AS=2.24e-14 PD=6e-07 PS=6e-07 $X=67640 $Y=59015 $D=0
M762 VDD 275 451 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=1.84e-14 AS=2.24e-14 PD=5.5e-07 PS=6e-07 $X=68020 $Y=55935 $D=0
M763 VDD 275 452 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=1.84e-14 AS=2.24e-14 PD=5.5e-07 PS=6e-07 $X=68020 $Y=59015 $D=0
M764 57 45 36 291 PMOS_VTL L=5e-08 W=1.6e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 $X=68075 $Y=50125 $D=0
M765 VDD 284 275 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 $X=68565 $Y=61790 $D=0
M766 VDD 55 284 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 $X=68575 $Y=62975 $D=0
M767 VDD 55 54 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 $X=68575 $Y=63835 $D=0
M768 55 54 58 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=2.4e-14 AS=1.92e-14 PD=6.2e-07 PS=5.6e-07 $X=68575 $Y=64695 $D=0
M769 58 52 55 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=2.4e-14 AS=2.4e-14 PD=6.2e-07 PS=6.2e-07 $X=68575 $Y=65095 $D=0
M770 VDD 50 58 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=1.92e-14 AS=2.4e-14 PD=5.6e-07 PS=6.2e-07 $X=68575 $Y=65495 $D=0
M771 VDD RESET 52 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 $X=68575 $Y=66355 $D=0
M772 VDD 51 50 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 $X=68575 $Y=67215 $D=0
M773 VDD 18 51 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 $X=68575 $Y=68075 $D=0
M774 56 51 55 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 $X=68575 $Y=68935 $D=0
M775 453 51 VDD VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=2.24e-14 AS=1.92e-14 PD=6e-07 PS=5.6e-07 $X=68575 $Y=69795 $D=0
M776 53 56 453 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=1.92e-14 AS=2.24e-14 PD=5.6e-07 PS=6e-07 $X=68575 $Y=70175 $D=0
M777 56 52 VDD VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=2.4e-14 AS=1.92e-14 PD=6.2e-07 PS=5.6e-07 $X=68575 $Y=71035 $D=0
M778 VDD 53 56 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=1.92e-14 AS=2.4e-14 PD=5.6e-07 PS=6.2e-07 $X=68575 $Y=71435 $D=0
M779 285 50 53 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 $X=68575 $Y=72295 $D=0
M780 VDD 286 285 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 $X=68575 $Y=73155 $D=0
M781 VDD B1 286 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 $X=68575 $Y=74015 $D=0
M782 454 45 291 291 PMOS_VTL L=5e-08 W=1.6e-07 AD=2.24e-14 AS=1.92e-14 PD=6e-07 PS=5.6e-07 $X=68935 $Y=50125 $D=0
M783 288 GND VDD VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=1.84e-14 AS=1.84e-14 PD=5.5e-07 PS=5.5e-07 $X=69150 $Y=56475 $D=0
M784 59 57 454 291 PMOS_VTL L=5e-08 W=1.6e-07 AD=1.92e-14 AS=2.24e-14 PD=5.6e-07 PS=6e-07 $X=69315 $Y=50125 $D=0
M785 61 GND 60 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=2.24e-14 AS=1.84e-14 PD=6e-07 PS=5.5e-07 $X=69920 $Y=56475 $D=0
M786 57 47 291 291 PMOS_VTL L=5e-08 W=1.6e-07 AD=2.4e-14 AS=1.92e-14 PD=6.2e-07 PS=5.6e-07 $X=70175 $Y=50125 $D=0
M787 62 288 61 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=1.84e-14 AS=2.24e-14 PD=5.5e-07 PS=6e-07 $X=70300 $Y=56475 $D=0
M788 291 59 57 291 PMOS_VTL L=5e-08 W=1.6e-07 AD=1.92e-14 AS=2.4e-14 PD=5.6e-07 PS=6.2e-07 $X=70575 $Y=50125 $D=0
M789 289 46 59 291 PMOS_VTL L=5e-08 W=1.6e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 $X=71435 $Y=50125 $D=0
M790 291 290 289 291 PMOS_VTL L=5e-08 W=1.6e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 $X=72295 $Y=50125 $D=0
M791 291 61 290 291 PMOS_VTL L=5e-08 W=1.6e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 $X=73155 $Y=50125 $D=0
M792 291 67 S2 291 PMOS_VTL L=5e-08 W=1.6e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 $X=74310 $Y=50125 $D=0
M793 VDD VDD 297 VDD PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=2.07e-14 PD=6.4e-07 PS=5.9e-07 $X=74590 $Y=55935 $D=0
M794 VDD VDD 299 VDD PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=2.07e-14 PD=6.4e-07 PS=5.9e-07 $X=74590 $Y=59015 $D=0
M795 VDD 69 VDD VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 $X=74950 $Y=62980 $D=0
M796 VDD 69 68 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 $X=74950 $Y=63840 $D=0
M797 69 68 72 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=2.4e-14 AS=1.92e-14 PD=6.2e-07 PS=5.6e-07 $X=74950 $Y=64700 $D=0
M798 72 65 69 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=2.4e-14 AS=2.4e-14 PD=6.2e-07 PS=6.2e-07 $X=74950 $Y=65100 $D=0
M799 VDD 63 72 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=1.92e-14 AS=2.4e-14 PD=5.6e-07 PS=6.2e-07 $X=74950 $Y=65500 $D=0
M800 VDD RESET 65 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 $X=74950 $Y=66360 $D=0
M801 VDD 64 63 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 $X=74950 $Y=67220 $D=0
M802 VDD 18 64 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 $X=74950 $Y=68080 $D=0
M803 70 64 69 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 $X=74950 $Y=68940 $D=0
M804 455 64 VDD VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=2.24e-14 AS=1.92e-14 PD=6e-07 PS=5.6e-07 $X=74950 $Y=69800 $D=0
M805 66 70 455 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=1.92e-14 AS=2.24e-14 PD=5.6e-07 PS=6e-07 $X=74950 $Y=70180 $D=0
M806 70 65 VDD VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=2.4e-14 AS=1.92e-14 PD=6.2e-07 PS=5.6e-07 $X=74950 $Y=71040 $D=0
M807 VDD 66 70 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=1.92e-14 AS=2.4e-14 PD=5.6e-07 PS=6.2e-07 $X=74950 $Y=71440 $D=0
M808 293 63 66 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 $X=74950 $Y=72300 $D=0
M809 VDD 294 293 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 $X=74950 $Y=73160 $D=0
M810 VDD A2 294 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 $X=74950 $Y=74020 $D=0
M811 297 295 VDD VDD PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=2.52e-14 PD=6.4e-07 PS=6.4e-07 $X=74970 $Y=55935 $D=0
M812 299 295 VDD VDD PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=2.52e-14 PD=6.4e-07 PS=6.4e-07 $X=74970 $Y=59015 $D=0
M813 291 67 71 291 PMOS_VTL L=5e-08 W=1.6e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 $X=75170 $Y=50125 $D=0
M814 77 48 297 VDD PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=2.52e-14 PD=6.4e-07 PS=6.4e-07 $X=75350 $Y=55935 $D=0
M815 78 49 299 VDD PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=2.52e-14 PD=6.4e-07 PS=6.4e-07 $X=75350 $Y=59015 $D=0
M816 456 VDD 77 VDD PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=2.52e-14 PD=6.4e-07 PS=6.4e-07 $X=75730 $Y=55935 $D=0
M817 457 VDD 78 VDD PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=2.52e-14 PD=6.4e-07 PS=6.4e-07 $X=75730 $Y=59015 $D=0
M818 67 71 73 291 PMOS_VTL L=5e-08 W=1.6e-07 AD=2.4e-14 AS=1.92e-14 PD=6.2e-07 PS=5.6e-07 $X=76030 $Y=50125 $D=0
M819 VDD 295 456 VDD PMOS_VTL L=5e-08 W=1.8e-07 AD=2.07e-14 AS=2.52e-14 PD=5.9e-07 PS=6.4e-07 $X=76110 $Y=55935 $D=0
M820 VDD 295 457 VDD PMOS_VTL L=5e-08 W=1.8e-07 AD=2.07e-14 AS=2.52e-14 PD=5.9e-07 PS=6.4e-07 $X=76110 $Y=59015 $D=0
M821 73 76 67 291 PMOS_VTL L=5e-08 W=1.6e-07 AD=2.4e-14 AS=2.4e-14 PD=6.2e-07 PS=6.2e-07 $X=76430 $Y=50125 $D=0
M822 291 75 73 291 PMOS_VTL L=5e-08 W=1.6e-07 AD=1.92e-14 AS=2.4e-14 PD=5.6e-07 PS=6.2e-07 $X=76830 $Y=50125 $D=0
M823 302 VDD VDD VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=2.24e-14 AS=1.84e-14 PD=6e-07 PS=5.5e-07 $X=76830 $Y=55935 $D=0
M824 304 VDD VDD VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=2.24e-14 AS=1.84e-14 PD=6e-07 PS=5.5e-07 $X=76830 $Y=59015 $D=0
M825 VDD 295 302 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=2.24e-14 AS=2.24e-14 PD=6e-07 PS=6e-07 $X=77210 $Y=55935 $D=0
M826 VDD 295 304 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=2.24e-14 AS=2.24e-14 PD=6e-07 PS=6e-07 $X=77210 $Y=59015 $D=0
M827 302 48 VDD VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=1.84e-14 AS=2.24e-14 PD=5.5e-07 PS=6e-07 $X=77590 $Y=55935 $D=0
M828 304 49 VDD VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=1.84e-14 AS=2.24e-14 PD=5.5e-07 PS=6e-07 $X=77590 $Y=59015 $D=0
M829 291 RESET 76 291 PMOS_VTL L=5e-08 W=1.6e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 $X=77690 $Y=50125 $D=0
M830 305 77 302 VDD PMOS_VTL L=5e-08 W=1.4e-07 AD=1.68e-14 AS=1.75e-14 PD=5.2e-07 PS=5.3e-07 $X=78330 $Y=55935 $D=0
M831 306 78 304 VDD PMOS_VTL L=5e-08 W=1.4e-07 AD=1.68e-14 AS=1.75e-14 PD=5.2e-07 PS=5.3e-07 $X=78330 $Y=59015 $D=0
M832 291 74 75 291 PMOS_VTL L=5e-08 W=1.6e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 $X=78550 $Y=50125 $D=0
M833 458 48 305 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=2.24e-14 AS=1.84e-14 PD=6e-07 PS=5.5e-07 $X=79060 $Y=55935 $D=0
M834 459 49 306 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=2.24e-14 AS=1.84e-14 PD=6e-07 PS=5.5e-07 $X=79060 $Y=59015 $D=0
M835 291 18 74 291 PMOS_VTL L=5e-08 W=1.6e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 $X=79410 $Y=50125 $D=0
M836 460 VDD 458 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=2.24e-14 AS=2.24e-14 PD=6e-07 PS=6e-07 $X=79440 $Y=55935 $D=0
M837 461 VDD 459 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=2.24e-14 AS=2.24e-14 PD=6e-07 PS=6e-07 $X=79440 $Y=59015 $D=0
M838 VDD 295 460 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=1.84e-14 AS=2.24e-14 PD=5.5e-07 PS=6e-07 $X=79820 $Y=55935 $D=0
M839 VDD 295 461 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=1.84e-14 AS=2.24e-14 PD=5.5e-07 PS=6e-07 $X=79820 $Y=59015 $D=0
M840 86 74 67 291 PMOS_VTL L=5e-08 W=1.6e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 $X=80270 $Y=50125 $D=0
M841 VDD 84 295 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 $X=80450 $Y=62980 $D=0
M842 VDD 84 83 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 $X=80450 $Y=63840 $D=0
M843 84 83 87 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=2.4e-14 AS=1.92e-14 PD=6.2e-07 PS=5.6e-07 $X=80450 $Y=64700 $D=0
M844 87 81 84 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=2.4e-14 AS=2.4e-14 PD=6.2e-07 PS=6.2e-07 $X=80450 $Y=65100 $D=0
M845 VDD 79 87 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=1.92e-14 AS=2.4e-14 PD=5.6e-07 PS=6.2e-07 $X=80450 $Y=65500 $D=0
M846 VDD RESET 81 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 $X=80450 $Y=66360 $D=0
M847 VDD 80 79 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 $X=80450 $Y=67220 $D=0
M848 VDD 18 80 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 $X=80450 $Y=68080 $D=0
M849 85 80 84 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 $X=80450 $Y=68940 $D=0
M850 462 80 VDD VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=2.24e-14 AS=1.92e-14 PD=6e-07 PS=5.6e-07 $X=80450 $Y=69800 $D=0
M851 82 85 462 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=1.92e-14 AS=2.24e-14 PD=5.6e-07 PS=6e-07 $X=80450 $Y=70180 $D=0
M852 85 81 VDD VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=2.4e-14 AS=1.92e-14 PD=6.2e-07 PS=5.6e-07 $X=80450 $Y=71040 $D=0
M853 VDD 82 85 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=1.92e-14 AS=2.4e-14 PD=5.6e-07 PS=6.2e-07 $X=80450 $Y=71440 $D=0
M854 307 79 82 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 $X=80450 $Y=72300 $D=0
M855 VDD 308 307 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 $X=80450 $Y=73160 $D=0
M856 VDD B2 308 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 $X=80450 $Y=74020 $D=0
M857 VDD 306 88 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 $X=80920 $Y=58615 $D=0
M858 310 GND VDD VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=1.84e-14 AS=1.84e-14 PD=5.5e-07 PS=5.5e-07 $X=80950 $Y=56475 $D=0
M859 463 74 291 291 PMOS_VTL L=5e-08 W=1.6e-07 AD=2.24e-14 AS=1.92e-14 PD=6e-07 PS=5.6e-07 $X=81130 $Y=50125 $D=0
M860 89 86 463 291 PMOS_VTL L=5e-08 W=1.6e-07 AD=1.92e-14 AS=2.24e-14 PD=5.6e-07 PS=6e-07 $X=81510 $Y=50125 $D=0
M861 90 GND 88 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=2.24e-14 AS=1.84e-14 PD=6e-07 PS=5.5e-07 $X=81720 $Y=56475 $D=0
M862 91 305 VDD VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 $X=81815 $Y=55295 $D=0
M863 91 310 90 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=1.84e-14 AS=2.24e-14 PD=5.5e-07 PS=6e-07 $X=82100 $Y=56475 $D=0
M864 86 76 291 291 PMOS_VTL L=5e-08 W=1.6e-07 AD=2.4e-14 AS=1.92e-14 PD=6.2e-07 PS=5.6e-07 $X=82370 $Y=50125 $D=0
M865 291 89 86 291 PMOS_VTL L=5e-08 W=1.6e-07 AD=1.92e-14 AS=2.4e-14 PD=5.6e-07 PS=6.2e-07 $X=82770 $Y=50125 $D=0
M866 311 75 89 291 PMOS_VTL L=5e-08 W=1.6e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 $X=83630 $Y=50125 $D=0
M867 291 312 311 291 PMOS_VTL L=5e-08 W=1.6e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 $X=84490 $Y=50125 $D=0
M868 291 90 312 291 PMOS_VTL L=5e-08 W=1.6e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 $X=85350 $Y=50125 $D=0
M869 VDD 313 320 VDD PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=2.07e-14 PD=6.4e-07 PS=5.9e-07 $X=86390 $Y=55775 $D=0
M870 VDD 313 322 VDD PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=2.07e-14 PD=6.4e-07 PS=5.9e-07 $X=86390 $Y=58855 $D=0
M871 336 99 S3 336 PMOS_VTL L=5e-08 W=1.6e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 $X=86575 $Y=50125 $D=0
M872 VDD 315 313 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 $X=86645 $Y=61795 $D=0
M873 VDD 97 315 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 $X=86655 $Y=62980 $D=0
M874 VDD 97 96 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 $X=86655 $Y=63840 $D=0
M875 97 96 100 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=2.4e-14 AS=1.92e-14 PD=6.2e-07 PS=5.6e-07 $X=86655 $Y=64700 $D=0
M876 100 94 97 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=2.4e-14 AS=2.4e-14 PD=6.2e-07 PS=6.2e-07 $X=86655 $Y=65100 $D=0
M877 VDD 92 100 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=1.92e-14 AS=2.4e-14 PD=5.6e-07 PS=6.2e-07 $X=86655 $Y=65500 $D=0
M878 VDD RESET 94 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 $X=86655 $Y=66360 $D=0
M879 VDD 93 92 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 $X=86655 $Y=67220 $D=0
M880 VDD 18 93 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 $X=86655 $Y=68080 $D=0
M881 98 93 97 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 $X=86655 $Y=68940 $D=0
M882 464 93 VDD VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=2.24e-14 AS=1.92e-14 PD=6e-07 PS=5.6e-07 $X=86655 $Y=69800 $D=0
M883 95 98 464 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=1.92e-14 AS=2.24e-14 PD=5.6e-07 PS=6e-07 $X=86655 $Y=70180 $D=0
M884 98 94 VDD VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=2.4e-14 AS=1.92e-14 PD=6.2e-07 PS=5.6e-07 $X=86655 $Y=71040 $D=0
M885 VDD 95 98 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=1.92e-14 AS=2.4e-14 PD=5.6e-07 PS=6.2e-07 $X=86655 $Y=71440 $D=0
M886 316 92 95 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 $X=86655 $Y=72300 $D=0
M887 VDD 317 316 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 $X=86655 $Y=73160 $D=0
M888 VDD A3 317 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 $X=86655 $Y=74020 $D=0
M889 320 318 VDD VDD PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=2.52e-14 PD=6.4e-07 PS=6.4e-07 $X=86770 $Y=55775 $D=0
M890 322 318 VDD VDD PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=2.52e-14 PD=6.4e-07 PS=6.4e-07 $X=86770 $Y=58855 $D=0
M891 106 77 320 VDD PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=2.52e-14 PD=6.4e-07 PS=6.4e-07 $X=87150 $Y=55775 $D=0
M892 107 78 322 VDD PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=2.52e-14 PD=6.4e-07 PS=6.4e-07 $X=87150 $Y=58855 $D=0
M893 336 99 101 336 PMOS_VTL L=5e-08 W=1.6e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 $X=87435 $Y=50125 $D=0
M894 465 313 106 VDD PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=2.52e-14 PD=6.4e-07 PS=6.4e-07 $X=87530 $Y=55775 $D=0
M895 466 313 107 VDD PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=2.52e-14 PD=6.4e-07 PS=6.4e-07 $X=87530 $Y=58855 $D=0
M896 VDD 318 465 VDD PMOS_VTL L=5e-08 W=1.8e-07 AD=2.07e-14 AS=2.52e-14 PD=5.9e-07 PS=6.4e-07 $X=87910 $Y=55775 $D=0
M897 VDD 318 466 VDD PMOS_VTL L=5e-08 W=1.8e-07 AD=2.07e-14 AS=2.52e-14 PD=5.9e-07 PS=6.4e-07 $X=87910 $Y=58855 $D=0
M898 99 101 102 336 PMOS_VTL L=5e-08 W=1.6e-07 AD=2.4e-14 AS=1.92e-14 PD=6.2e-07 PS=5.6e-07 $X=88295 $Y=50125 $D=0
M899 325 313 VDD VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=2.24e-14 AS=1.84e-14 PD=6e-07 PS=5.5e-07 $X=88630 $Y=55775 $D=0
M900 327 313 VDD VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=2.24e-14 AS=1.84e-14 PD=6e-07 PS=5.5e-07 $X=88630 $Y=58855 $D=0
M901 102 105 99 336 PMOS_VTL L=5e-08 W=1.6e-07 AD=2.4e-14 AS=2.4e-14 PD=6.2e-07 PS=6.2e-07 $X=88695 $Y=50125 $D=0
M902 VDD 318 325 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=2.24e-14 AS=2.24e-14 PD=6e-07 PS=6e-07 $X=89010 $Y=55775 $D=0
M903 VDD 318 327 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=2.24e-14 AS=2.24e-14 PD=6e-07 PS=6e-07 $X=89010 $Y=58855 $D=0
M904 336 104 102 336 PMOS_VTL L=5e-08 W=1.6e-07 AD=1.92e-14 AS=2.4e-14 PD=5.6e-07 PS=6.2e-07 $X=89095 $Y=50125 $D=0
M905 325 77 VDD VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=1.84e-14 AS=2.24e-14 PD=5.5e-07 PS=6e-07 $X=89390 $Y=55775 $D=0
M906 327 78 VDD VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=1.84e-14 AS=2.24e-14 PD=5.5e-07 PS=6e-07 $X=89390 $Y=58855 $D=0
M907 336 RESET 105 336 PMOS_VTL L=5e-08 W=1.6e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 $X=89955 $Y=50125 $D=0
M908 120 106 325 VDD PMOS_VTL L=5e-08 W=1.4e-07 AD=1.68e-14 AS=1.75e-14 PD=5.2e-07 PS=5.3e-07 $X=90130 $Y=55775 $D=0
M909 117 107 327 VDD PMOS_VTL L=5e-08 W=1.4e-07 AD=1.68e-14 AS=1.75e-14 PD=5.2e-07 PS=5.3e-07 $X=90130 $Y=58855 $D=0
M910 336 103 104 336 PMOS_VTL L=5e-08 W=1.6e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 $X=90815 $Y=50125 $D=0
M911 467 77 120 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=2.24e-14 AS=1.84e-14 PD=6e-07 PS=5.5e-07 $X=90860 $Y=55775 $D=0
M912 468 78 117 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=2.24e-14 AS=1.84e-14 PD=6e-07 PS=5.5e-07 $X=90860 $Y=58855 $D=0
M913 469 313 467 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=2.24e-14 AS=2.24e-14 PD=6e-07 PS=6e-07 $X=91240 $Y=55775 $D=0
M914 470 313 468 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=2.24e-14 AS=2.24e-14 PD=6e-07 PS=6e-07 $X=91240 $Y=58855 $D=0
M915 VDD 318 469 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=1.84e-14 AS=2.24e-14 PD=5.5e-07 PS=6e-07 $X=91620 $Y=55775 $D=0
M916 VDD 318 470 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=1.84e-14 AS=2.24e-14 PD=5.5e-07 PS=6e-07 $X=91620 $Y=58855 $D=0
M917 336 18 103 336 PMOS_VTL L=5e-08 W=1.6e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 $X=91675 $Y=50125 $D=0
M918 VDD 328 318 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 $X=92165 $Y=61795 $D=0
M919 VDD 113 328 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 $X=92175 $Y=62980 $D=0
M920 VDD 113 112 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 $X=92175 $Y=63840 $D=0
M921 113 112 115 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=2.4e-14 AS=1.92e-14 PD=6.2e-07 PS=5.6e-07 $X=92175 $Y=64700 $D=0
M922 115 110 113 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=2.4e-14 AS=2.4e-14 PD=6.2e-07 PS=6.2e-07 $X=92175 $Y=65100 $D=0
M923 VDD 108 115 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=1.92e-14 AS=2.4e-14 PD=5.6e-07 PS=6.2e-07 $X=92175 $Y=65500 $D=0
M924 VDD RESET 110 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 $X=92175 $Y=66360 $D=0
M925 VDD 109 108 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 $X=92175 $Y=67220 $D=0
M926 VDD 18 109 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 $X=92175 $Y=68080 $D=0
M927 114 109 113 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 $X=92175 $Y=68940 $D=0
M928 471 109 VDD VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=2.24e-14 AS=1.92e-14 PD=6e-07 PS=5.6e-07 $X=92175 $Y=69800 $D=0
M929 111 114 471 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=1.92e-14 AS=2.24e-14 PD=5.6e-07 PS=6e-07 $X=92175 $Y=70180 $D=0
M930 114 110 VDD VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=2.4e-14 AS=1.92e-14 PD=6.2e-07 PS=5.6e-07 $X=92175 $Y=71040 $D=0
M931 VDD 111 114 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=1.92e-14 AS=2.4e-14 PD=5.6e-07 PS=6.2e-07 $X=92175 $Y=71440 $D=0
M932 329 108 111 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 $X=92175 $Y=72300 $D=0
M933 VDD 330 329 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 $X=92175 $Y=73160 $D=0
M934 VDD B3 330 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 $X=92175 $Y=74020 $D=0
M935 116 103 99 336 PMOS_VTL L=5e-08 W=1.6e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 $X=92535 $Y=50125 $D=0
M936 332 GND VDD VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=1.84e-14 AS=1.84e-14 PD=5.5e-07 PS=5.5e-07 $X=92750 $Y=56315 $D=0
M937 472 103 336 336 PMOS_VTL L=5e-08 W=1.6e-07 AD=2.24e-14 AS=1.92e-14 PD=6e-07 PS=5.6e-07 $X=93395 $Y=50125 $D=0
M938 118 GND 117 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=2.24e-14 AS=1.84e-14 PD=6e-07 PS=5.5e-07 $X=93520 $Y=56315 $D=0
M939 119 116 472 336 PMOS_VTL L=5e-08 W=1.6e-07 AD=1.92e-14 AS=2.24e-14 PD=5.6e-07 PS=6e-07 $X=93775 $Y=50125 $D=0
M940 120 332 118 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=1.84e-14 AS=2.24e-14 PD=5.5e-07 PS=6e-07 $X=93900 $Y=56315 $D=0
M941 116 105 336 336 PMOS_VTL L=5e-08 W=1.6e-07 AD=2.4e-14 AS=1.92e-14 PD=6.2e-07 PS=5.6e-07 $X=94635 $Y=50125 $D=0
M942 336 119 116 336 PMOS_VTL L=5e-08 W=1.6e-07 AD=1.92e-14 AS=2.4e-14 PD=5.6e-07 PS=6.2e-07 $X=95035 $Y=50125 $D=0
M943 333 GND VDD VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=1.84e-14 AS=1.84e-14 PD=5.5e-07 PS=5.5e-07 $X=95855 $Y=56290 $D=0
M944 334 104 119 336 PMOS_VTL L=5e-08 W=1.6e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 $X=95895 $Y=50125 $D=0
M945 121 GND 107 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=2.24e-14 AS=1.84e-14 PD=6e-07 PS=5.5e-07 $X=96625 $Y=56290 $D=0
M946 336 335 334 336 PMOS_VTL L=5e-08 W=1.6e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 $X=96755 $Y=50125 $D=0
M947 106 333 121 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=1.84e-14 AS=2.24e-14 PD=5.5e-07 PS=6e-07 $X=97005 $Y=56290 $D=0
M948 336 118 335 336 PMOS_VTL L=5e-08 W=1.6e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 $X=97615 $Y=50125 $D=0
M949 359 122 S4 359 PMOS_VTL L=5e-08 W=1.6e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 $X=99550 $Y=50125 $D=0
M950 359 122 123 359 PMOS_VTL L=5e-08 W=1.6e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 $X=100410 $Y=50125 $D=0
M951 122 123 126 359 PMOS_VTL L=5e-08 W=1.6e-07 AD=2.4e-14 AS=1.92e-14 PD=6.2e-07 PS=5.6e-07 $X=101270 $Y=50125 $D=0
M952 147 338 343 147 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=2.07e-14 PD=6.4e-07 PS=5.9e-07 $X=101460 $Y=55935 $D=0
M953 VDD 338 345 VDD PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=2.07e-14 PD=6.4e-07 PS=5.9e-07 $X=101460 $Y=58855 $D=0
M954 126 135 122 359 PMOS_VTL L=5e-08 W=1.6e-07 AD=2.4e-14 AS=2.4e-14 PD=6.2e-07 PS=6.2e-07 $X=101670 $Y=50125 $D=0
M955 VDD 130 338 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 $X=101820 $Y=62980 $D=0
M956 VDD 130 129 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 $X=101820 $Y=63840 $D=0
M957 130 129 132 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=2.4e-14 AS=1.92e-14 PD=6.2e-07 PS=5.6e-07 $X=101820 $Y=64700 $D=0
M958 132 127 130 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=2.4e-14 AS=2.4e-14 PD=6.2e-07 PS=6.2e-07 $X=101820 $Y=65100 $D=0
M959 VDD 124 132 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=1.92e-14 AS=2.4e-14 PD=5.6e-07 PS=6.2e-07 $X=101820 $Y=65500 $D=0
M960 VDD RESET 127 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 $X=101820 $Y=66360 $D=0
M961 VDD 125 124 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 $X=101820 $Y=67220 $D=0
M962 VDD 18 125 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 $X=101820 $Y=68080 $D=0
M963 131 125 130 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 $X=101820 $Y=68940 $D=0
M964 473 125 VDD VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=2.24e-14 AS=1.92e-14 PD=6e-07 PS=5.6e-07 $X=101820 $Y=69800 $D=0
M965 128 131 473 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=1.92e-14 AS=2.24e-14 PD=5.6e-07 PS=6e-07 $X=101820 $Y=70180 $D=0
M966 131 127 VDD VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=2.4e-14 AS=1.92e-14 PD=6.2e-07 PS=5.6e-07 $X=101820 $Y=71040 $D=0
M967 VDD 128 131 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=1.92e-14 AS=2.4e-14 PD=5.6e-07 PS=6.2e-07 $X=101820 $Y=71440 $D=0
M968 339 124 128 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 $X=101820 $Y=72300 $D=0
M969 VDD 340 339 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 $X=101820 $Y=73160 $D=0
M970 VDD A4 340 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 $X=101820 $Y=74020 $D=0
M971 343 341 147 147 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=2.52e-14 PD=6.4e-07 PS=6.4e-07 $X=101840 $Y=55935 $D=0
M972 345 341 VDD VDD PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=2.52e-14 PD=6.4e-07 PS=6.4e-07 $X=101840 $Y=58855 $D=0
M973 359 134 126 359 PMOS_VTL L=5e-08 W=1.6e-07 AD=1.92e-14 AS=2.4e-14 PD=5.6e-07 PS=6.2e-07 $X=102070 $Y=50125 $D=0
M974 136 147 343 147 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=2.52e-14 PD=6.4e-07 PS=6.4e-07 $X=102220 $Y=55935 $D=0
M975 137 GND 345 VDD PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=2.52e-14 PD=6.4e-07 PS=6.4e-07 $X=102220 $Y=58855 $D=0
M976 474 338 136 147 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=2.52e-14 PD=6.4e-07 PS=6.4e-07 $X=102600 $Y=55935 $D=0
M977 475 338 137 VDD PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=2.52e-14 PD=6.4e-07 PS=6.4e-07 $X=102600 $Y=58855 $D=0
M978 359 RESET 135 359 PMOS_VTL L=5e-08 W=1.6e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 $X=102930 $Y=50125 $D=0
M979 147 341 474 147 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.07e-14 AS=2.52e-14 PD=5.9e-07 PS=6.4e-07 $X=102980 $Y=55935 $D=0
M980 VDD 341 475 VDD PMOS_VTL L=5e-08 W=1.8e-07 AD=2.07e-14 AS=2.52e-14 PD=5.9e-07 PS=6.4e-07 $X=102980 $Y=58855 $D=0
M981 348 338 147 147 PMOS_VTL L=5e-08 W=1.6e-07 AD=2.24e-14 AS=1.84e-14 PD=6e-07 PS=5.5e-07 $X=103700 $Y=55935 $D=0
M982 350 338 VDD VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=2.24e-14 AS=1.84e-14 PD=6e-07 PS=5.5e-07 $X=103700 $Y=58855 $D=0
M983 359 133 134 359 PMOS_VTL L=5e-08 W=1.6e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 $X=103790 $Y=50125 $D=0
M984 147 341 348 147 PMOS_VTL L=5e-08 W=1.6e-07 AD=2.24e-14 AS=2.24e-14 PD=6e-07 PS=6e-07 $X=104080 $Y=55935 $D=0
M985 VDD 341 350 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=2.24e-14 AS=2.24e-14 PD=6e-07 PS=6e-07 $X=104080 $Y=58855 $D=0
M986 348 147 147 147 PMOS_VTL L=5e-08 W=1.6e-07 AD=1.84e-14 AS=2.24e-14 PD=5.5e-07 PS=6e-07 $X=104460 $Y=55935 $D=0
M987 350 GND VDD VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=1.84e-14 AS=2.24e-14 PD=5.5e-07 PS=6e-07 $X=104460 $Y=58855 $D=0
M988 359 18 133 359 PMOS_VTL L=5e-08 W=1.6e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 $X=104650 $Y=50125 $D=0
M989 351 136 348 147 PMOS_VTL L=5e-08 W=1.4e-07 AD=1.68e-14 AS=1.75e-14 PD=5.2e-07 PS=5.3e-07 $X=105200 $Y=55935 $D=0
M990 352 137 350 VDD PMOS_VTL L=5e-08 W=1.4e-07 AD=1.68e-14 AS=1.75e-14 PD=5.2e-07 PS=5.3e-07 $X=105200 $Y=58855 $D=0
M991 139 133 122 359 PMOS_VTL L=5e-08 W=1.6e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 $X=105510 $Y=50125 $D=0
M992 476 147 351 147 PMOS_VTL L=5e-08 W=1.6e-07 AD=2.24e-14 AS=1.84e-14 PD=6e-07 PS=5.5e-07 $X=105930 $Y=55935 $D=0
M993 477 GND 352 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=2.24e-14 AS=1.84e-14 PD=6e-07 PS=5.5e-07 $X=105930 $Y=58855 $D=0
M994 478 338 476 147 PMOS_VTL L=5e-08 W=1.6e-07 AD=2.24e-14 AS=2.24e-14 PD=6e-07 PS=6e-07 $X=106310 $Y=55935 $D=0
M995 479 338 477 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=2.24e-14 AS=2.24e-14 PD=6e-07 PS=6e-07 $X=106310 $Y=58855 $D=0
M996 480 133 359 359 PMOS_VTL L=5e-08 W=1.6e-07 AD=2.24e-14 AS=1.92e-14 PD=6e-07 PS=5.6e-07 $X=106370 $Y=50125 $D=0
M997 147 341 478 147 PMOS_VTL L=5e-08 W=1.6e-07 AD=1.84e-14 AS=2.24e-14 PD=5.5e-07 PS=6e-07 $X=106690 $Y=55935 $D=0
M998 VDD 341 479 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=1.84e-14 AS=2.24e-14 PD=5.5e-07 PS=6e-07 $X=106690 $Y=58855 $D=0
M999 146 139 480 359 PMOS_VTL L=5e-08 W=1.6e-07 AD=1.92e-14 AS=2.24e-14 PD=5.6e-07 PS=6e-07 $X=106750 $Y=50125 $D=0
M1000 VDD 144 341 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 $X=107320 $Y=62980 $D=0
M1001 VDD 144 143 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 $X=107320 $Y=63840 $D=0
M1002 144 143 148 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=2.4e-14 AS=1.92e-14 PD=6.2e-07 PS=5.6e-07 $X=107320 $Y=64700 $D=0
M1003 148 141 144 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=2.4e-14 AS=2.4e-14 PD=6.2e-07 PS=6.2e-07 $X=107320 $Y=65100 $D=0
M1004 VDD 138 148 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=1.92e-14 AS=2.4e-14 PD=5.6e-07 PS=6.2e-07 $X=107320 $Y=65500 $D=0
M1005 VDD RESET 141 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 $X=107320 $Y=66360 $D=0
M1006 VDD 140 138 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 $X=107320 $Y=67220 $D=0
M1007 VDD 18 140 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 $X=107320 $Y=68080 $D=0
M1008 145 140 144 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 $X=107320 $Y=68940 $D=0
M1009 481 140 VDD VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=2.24e-14 AS=1.92e-14 PD=6e-07 PS=5.6e-07 $X=107320 $Y=69800 $D=0
M1010 142 145 481 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=1.92e-14 AS=2.24e-14 PD=5.6e-07 PS=6e-07 $X=107320 $Y=70180 $D=0
M1011 145 141 VDD VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=2.4e-14 AS=1.92e-14 PD=6.2e-07 PS=5.6e-07 $X=107320 $Y=71040 $D=0
M1012 VDD 142 145 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=1.92e-14 AS=2.4e-14 PD=5.6e-07 PS=6.2e-07 $X=107320 $Y=71440 $D=0
M1013 353 138 142 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 $X=107320 $Y=72300 $D=0
M1014 VDD 354 353 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 $X=107320 $Y=73160 $D=0
M1015 VDD B4 354 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 $X=107320 $Y=74020 $D=0
M1016 139 135 359 359 PMOS_VTL L=5e-08 W=1.6e-07 AD=2.4e-14 AS=1.92e-14 PD=6.2e-07 PS=5.6e-07 $X=107610 $Y=50125 $D=0
M1017 VDD 352 149 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 $X=107790 $Y=58455 $D=0
M1018 356 121 147 147 PMOS_VTL L=5e-08 W=1.6e-07 AD=1.84e-14 AS=1.84e-14 PD=5.5e-07 PS=5.5e-07 $X=107820 $Y=56315 $D=0
M1019 359 146 139 359 PMOS_VTL L=5e-08 W=1.6e-07 AD=1.92e-14 AS=2.4e-14 PD=5.6e-07 PS=6.2e-07 $X=108010 $Y=50125 $D=0
M1020 150 121 149 147 PMOS_VTL L=5e-08 W=1.6e-07 AD=2.24e-14 AS=1.84e-14 PD=6e-07 PS=5.5e-07 $X=108590 $Y=56315 $D=0
M1021 151 351 147 147 PMOS_VTL L=5e-08 W=1.6e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 $X=108685 $Y=55295 $D=0
M1022 357 134 146 359 PMOS_VTL L=5e-08 W=1.6e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 $X=108870 $Y=50125 $D=0
M1023 151 356 150 147 PMOS_VTL L=5e-08 W=1.6e-07 AD=1.84e-14 AS=2.24e-14 PD=5.5e-07 PS=6e-07 $X=108970 $Y=56315 $D=0
M1024 359 358 357 359 PMOS_VTL L=5e-08 W=1.6e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 $X=109730 $Y=50125 $D=0
M1025 359 150 358 359 PMOS_VTL L=5e-08 W=1.6e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 $X=110590 $Y=50125 $D=0
M1026 384 154 S5 384 PMOS_VTL L=5e-08 W=1.6e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 $X=111970 $Y=50125 $D=0
M1027 384 154 155 384 PMOS_VTL L=5e-08 W=1.6e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 $X=112830 $Y=50125 $D=0
M1028 379 361 367 379 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=2.07e-14 PD=6.4e-07 PS=5.9e-07 $X=113260 $Y=55725 $D=0
M1029 VDD 361 369 VDD PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=2.07e-14 PD=6.4e-07 PS=5.9e-07 $X=113260 $Y=58805 $D=0
M1030 VDD 362 361 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 $X=113515 $Y=61795 $D=0
M1031 VDD 159 362 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 $X=113525 $Y=62980 $D=0
M1032 VDD 159 158 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 $X=113525 $Y=63840 $D=0
M1033 159 158 162 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=2.4e-14 AS=1.92e-14 PD=6.2e-07 PS=5.6e-07 $X=113525 $Y=64700 $D=0
M1034 162 156 159 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=2.4e-14 AS=2.4e-14 PD=6.2e-07 PS=6.2e-07 $X=113525 $Y=65100 $D=0
M1035 VDD 152 162 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=1.92e-14 AS=2.4e-14 PD=5.6e-07 PS=6.2e-07 $X=113525 $Y=65500 $D=0
M1036 VDD RESET 156 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 $X=113525 $Y=66360 $D=0
M1037 VDD 153 152 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 $X=113525 $Y=67220 $D=0
M1038 VDD 18 153 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 $X=113525 $Y=68080 $D=0
M1039 160 153 159 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 $X=113525 $Y=68940 $D=0
M1040 482 153 VDD VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=2.24e-14 AS=1.92e-14 PD=6e-07 PS=5.6e-07 $X=113525 $Y=69800 $D=0
M1041 157 160 482 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=1.92e-14 AS=2.24e-14 PD=5.6e-07 PS=6e-07 $X=113525 $Y=70180 $D=0
M1042 160 156 VDD VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=2.4e-14 AS=1.92e-14 PD=6.2e-07 PS=5.6e-07 $X=113525 $Y=71040 $D=0
M1043 VDD 157 160 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=1.92e-14 AS=2.4e-14 PD=5.6e-07 PS=6.2e-07 $X=113525 $Y=71440 $D=0
M1044 363 152 157 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 $X=113525 $Y=72300 $D=0
M1045 VDD 364 363 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 $X=113525 $Y=73160 $D=0
M1046 VDD A5 364 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 $X=113525 $Y=74020 $D=0
M1047 367 365 379 379 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=2.52e-14 PD=6.4e-07 PS=6.4e-07 $X=113640 $Y=55725 $D=0
M1048 369 365 VDD VDD PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=2.52e-14 PD=6.4e-07 PS=6.4e-07 $X=113640 $Y=58805 $D=0
M1049 154 155 161 384 PMOS_VTL L=5e-08 W=1.6e-07 AD=2.4e-14 AS=1.92e-14 PD=6.2e-07 PS=5.6e-07 $X=113690 $Y=50125 $D=0
M1050 166 136 367 379 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=2.52e-14 PD=6.4e-07 PS=6.4e-07 $X=114020 $Y=55725 $D=0
M1051 167 137 369 VDD PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=2.52e-14 PD=6.4e-07 PS=6.4e-07 $X=114020 $Y=58805 $D=0
M1052 161 165 154 384 PMOS_VTL L=5e-08 W=1.6e-07 AD=2.4e-14 AS=2.4e-14 PD=6.2e-07 PS=6.2e-07 $X=114090 $Y=50125 $D=0
M1053 483 361 166 379 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=2.52e-14 PD=6.4e-07 PS=6.4e-07 $X=114400 $Y=55725 $D=0
M1054 484 361 167 VDD PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=2.52e-14 PD=6.4e-07 PS=6.4e-07 $X=114400 $Y=58805 $D=0
M1055 384 164 161 384 PMOS_VTL L=5e-08 W=1.6e-07 AD=1.92e-14 AS=2.4e-14 PD=5.6e-07 PS=6.2e-07 $X=114490 $Y=50125 $D=0
M1056 379 365 483 379 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.07e-14 AS=2.52e-14 PD=5.9e-07 PS=6.4e-07 $X=114780 $Y=55725 $D=0
M1057 VDD 365 484 VDD PMOS_VTL L=5e-08 W=1.8e-07 AD=2.07e-14 AS=2.52e-14 PD=5.9e-07 PS=6.4e-07 $X=114780 $Y=58805 $D=0
M1058 384 RESET 165 384 PMOS_VTL L=5e-08 W=1.6e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 $X=115350 $Y=50125 $D=0
M1059 372 361 379 379 PMOS_VTL L=5e-08 W=1.6e-07 AD=2.24e-14 AS=1.84e-14 PD=6e-07 PS=5.5e-07 $X=115500 $Y=55725 $D=0
M1060 374 361 VDD VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=2.24e-14 AS=1.84e-14 PD=6e-07 PS=5.5e-07 $X=115500 $Y=58805 $D=0
M1061 379 365 372 379 PMOS_VTL L=5e-08 W=1.6e-07 AD=2.24e-14 AS=2.24e-14 PD=6e-07 PS=6e-07 $X=115880 $Y=55725 $D=0
M1062 VDD 365 374 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=2.24e-14 AS=2.24e-14 PD=6e-07 PS=6e-07 $X=115880 $Y=58805 $D=0
M1063 384 163 164 384 PMOS_VTL L=5e-08 W=1.6e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 $X=116210 $Y=50125 $D=0
M1064 372 136 379 379 PMOS_VTL L=5e-08 W=1.6e-07 AD=1.84e-14 AS=2.24e-14 PD=5.5e-07 PS=6e-07 $X=116260 $Y=55725 $D=0
M1065 374 137 VDD VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=1.84e-14 AS=2.24e-14 PD=5.5e-07 PS=6e-07 $X=116260 $Y=58805 $D=0
M1066 375 166 372 379 PMOS_VTL L=5e-08 W=1.4e-07 AD=1.68e-14 AS=1.75e-14 PD=5.2e-07 PS=5.3e-07 $X=117000 $Y=55725 $D=0
M1067 178 167 374 VDD PMOS_VTL L=5e-08 W=1.4e-07 AD=1.68e-14 AS=1.75e-14 PD=5.2e-07 PS=5.3e-07 $X=117000 $Y=58805 $D=0
M1068 384 18 163 384 PMOS_VTL L=5e-08 W=1.6e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 $X=117070 $Y=50125 $D=0
M1069 485 136 375 379 PMOS_VTL L=5e-08 W=1.6e-07 AD=2.24e-14 AS=1.84e-14 PD=6e-07 PS=5.5e-07 $X=117730 $Y=55725 $D=0
M1070 486 137 178 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=2.24e-14 AS=1.84e-14 PD=6e-07 PS=5.5e-07 $X=117730 $Y=58805 $D=0
M1071 170 163 154 384 PMOS_VTL L=5e-08 W=1.6e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 $X=117930 $Y=50125 $D=0
M1072 487 361 485 379 PMOS_VTL L=5e-08 W=1.6e-07 AD=2.24e-14 AS=2.24e-14 PD=6e-07 PS=6e-07 $X=118110 $Y=55725 $D=0
M1073 488 361 486 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=2.24e-14 AS=2.24e-14 PD=6e-07 PS=6e-07 $X=118110 $Y=58805 $D=0
M1074 379 365 487 379 PMOS_VTL L=5e-08 W=1.6e-07 AD=1.84e-14 AS=2.24e-14 PD=5.5e-07 PS=6e-07 $X=118490 $Y=55725 $D=0
M1075 VDD 365 488 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=1.84e-14 AS=2.24e-14 PD=5.5e-07 PS=6e-07 $X=118490 $Y=58805 $D=0
M1076 489 163 384 384 PMOS_VTL L=5e-08 W=1.6e-07 AD=2.24e-14 AS=1.92e-14 PD=6e-07 PS=5.6e-07 $X=118790 $Y=50125 $D=0
M1077 VDD 376 365 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 $X=119035 $Y=61795 $D=0
M1078 VDD 174 376 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 $X=119045 $Y=62980 $D=0
M1079 VDD 174 173 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 $X=119045 $Y=63840 $D=0
M1080 174 173 176 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=2.4e-14 AS=1.92e-14 PD=6.2e-07 PS=5.6e-07 $X=119045 $Y=64700 $D=0
M1081 176 171 174 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=2.4e-14 AS=2.4e-14 PD=6.2e-07 PS=6.2e-07 $X=119045 $Y=65100 $D=0
M1082 VDD 168 176 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=1.92e-14 AS=2.4e-14 PD=5.6e-07 PS=6.2e-07 $X=119045 $Y=65500 $D=0
M1083 VDD RESET 171 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 $X=119045 $Y=66360 $D=0
M1084 VDD 169 168 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 $X=119045 $Y=67220 $D=0
M1085 VDD 18 169 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 $X=119045 $Y=68080 $D=0
M1086 175 169 174 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 $X=119045 $Y=68940 $D=0
M1087 490 169 VDD VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=2.24e-14 AS=1.92e-14 PD=6e-07 PS=5.6e-07 $X=119045 $Y=69800 $D=0
M1088 172 175 490 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=1.92e-14 AS=2.24e-14 PD=5.6e-07 PS=6e-07 $X=119045 $Y=70180 $D=0
M1089 175 171 VDD VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=2.4e-14 AS=1.92e-14 PD=6.2e-07 PS=5.6e-07 $X=119045 $Y=71040 $D=0
M1090 VDD 172 175 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=1.92e-14 AS=2.4e-14 PD=5.6e-07 PS=6.2e-07 $X=119045 $Y=71440 $D=0
M1091 377 168 172 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 $X=119045 $Y=72300 $D=0
M1092 VDD 378 377 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 $X=119045 $Y=73160 $D=0
M1093 VDD B5 378 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 $X=119045 $Y=74020 $D=0
M1094 177 170 489 384 PMOS_VTL L=5e-08 W=1.6e-07 AD=1.92e-14 AS=2.24e-14 PD=5.6e-07 PS=6e-07 $X=119170 $Y=50125 $D=0
M1095 381 121 379 379 PMOS_VTL L=5e-08 W=1.6e-07 AD=1.84e-14 AS=1.84e-14 PD=5.5e-07 PS=5.5e-07 $X=119620 $Y=56265 $D=0
M1096 170 165 384 384 PMOS_VTL L=5e-08 W=1.6e-07 AD=2.4e-14 AS=1.92e-14 PD=6.2e-07 PS=5.6e-07 $X=120030 $Y=50125 $D=0
M1097 179 121 178 379 PMOS_VTL L=5e-08 W=1.6e-07 AD=2.24e-14 AS=1.84e-14 PD=6e-07 PS=5.5e-07 $X=120390 $Y=56265 $D=0
M1098 384 177 170 384 PMOS_VTL L=5e-08 W=1.6e-07 AD=1.92e-14 AS=2.4e-14 PD=5.6e-07 PS=6.2e-07 $X=120430 $Y=50125 $D=0
M1099 180 381 179 379 PMOS_VTL L=5e-08 W=1.6e-07 AD=1.84e-14 AS=2.24e-14 PD=5.5e-07 PS=6e-07 $X=120770 $Y=56265 $D=0
M1100 382 164 177 384 PMOS_VTL L=5e-08 W=1.6e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 $X=121290 $Y=50125 $D=0
M1101 384 383 382 384 PMOS_VTL L=5e-08 W=1.6e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 $X=122150 $Y=50125 $D=0
M1102 384 179 383 384 PMOS_VTL L=5e-08 W=1.6e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 $X=123010 $Y=50125 $D=0
M1103 407 183 S6 407 PMOS_VTL L=5e-08 W=1.6e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 $X=124525 $Y=50125 $D=0
M1104 205 386 391 205 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=2.07e-14 PD=6.4e-07 PS=5.9e-07 $X=125060 $Y=55775 $D=0
M1105 VDD 386 393 VDD PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=2.07e-14 PD=6.4e-07 PS=5.9e-07 $X=125060 $Y=58855 $D=0
M1106 407 183 186 407 PMOS_VTL L=5e-08 W=1.6e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 $X=125385 $Y=50125 $D=0
M1107 VDD 188 386 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 $X=125420 $Y=62980 $D=0
M1108 VDD 188 187 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 $X=125420 $Y=63840 $D=0
M1109 188 187 190 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=2.4e-14 AS=1.92e-14 PD=6.2e-07 PS=5.6e-07 $X=125420 $Y=64700 $D=0
M1110 190 184 188 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=2.4e-14 AS=2.4e-14 PD=6.2e-07 PS=6.2e-07 $X=125420 $Y=65100 $D=0
M1111 VDD 181 190 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=1.92e-14 AS=2.4e-14 PD=5.6e-07 PS=6.2e-07 $X=125420 $Y=65500 $D=0
M1112 VDD RESET 184 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 $X=125420 $Y=66360 $D=0
M1113 VDD 182 181 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 $X=125420 $Y=67220 $D=0
M1114 VDD 18 182 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 $X=125420 $Y=68080 $D=0
M1115 189 182 188 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 $X=125420 $Y=68940 $D=0
M1116 491 182 VDD VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=2.24e-14 AS=1.92e-14 PD=6e-07 PS=5.6e-07 $X=125420 $Y=69800 $D=0
M1117 185 189 491 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=1.92e-14 AS=2.24e-14 PD=5.6e-07 PS=6e-07 $X=125420 $Y=70180 $D=0
M1118 189 184 VDD VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=2.4e-14 AS=1.92e-14 PD=6.2e-07 PS=5.6e-07 $X=125420 $Y=71040 $D=0
M1119 VDD 185 189 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=1.92e-14 AS=2.4e-14 PD=5.6e-07 PS=6.2e-07 $X=125420 $Y=71440 $D=0
M1120 387 181 185 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 $X=125420 $Y=72300 $D=0
M1121 VDD 388 387 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 $X=125420 $Y=73160 $D=0
M1122 VDD A6 388 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 $X=125420 $Y=74020 $D=0
M1123 391 389 205 205 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=2.52e-14 PD=6.4e-07 PS=6.4e-07 $X=125440 $Y=55775 $D=0
M1124 393 389 VDD VDD PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=2.52e-14 PD=6.4e-07 PS=6.4e-07 $X=125440 $Y=58855 $D=0
M1125 195 166 391 205 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=2.52e-14 PD=6.4e-07 PS=6.4e-07 $X=125820 $Y=55775 $D=0
M1126 196 167 393 VDD PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=2.52e-14 PD=6.4e-07 PS=6.4e-07 $X=125820 $Y=58855 $D=0
M1127 492 386 195 205 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=2.52e-14 PD=6.4e-07 PS=6.4e-07 $X=126200 $Y=55775 $D=0
M1128 493 386 196 VDD PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=2.52e-14 PD=6.4e-07 PS=6.4e-07 $X=126200 $Y=58855 $D=0
M1129 183 186 191 407 PMOS_VTL L=5e-08 W=1.6e-07 AD=2.4e-14 AS=1.92e-14 PD=6.2e-07 PS=5.6e-07 $X=126245 $Y=50125 $D=0
M1130 205 389 492 205 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.07e-14 AS=2.52e-14 PD=5.9e-07 PS=6.4e-07 $X=126580 $Y=55775 $D=0
M1131 VDD 389 493 VDD PMOS_VTL L=5e-08 W=1.8e-07 AD=2.07e-14 AS=2.52e-14 PD=5.9e-07 PS=6.4e-07 $X=126580 $Y=58855 $D=0
M1132 191 194 183 407 PMOS_VTL L=5e-08 W=1.6e-07 AD=2.4e-14 AS=2.4e-14 PD=6.2e-07 PS=6.2e-07 $X=126645 $Y=50125 $D=0
M1133 407 193 191 407 PMOS_VTL L=5e-08 W=1.6e-07 AD=1.92e-14 AS=2.4e-14 PD=5.6e-07 PS=6.2e-07 $X=127045 $Y=50125 $D=0
M1134 396 386 205 205 PMOS_VTL L=5e-08 W=1.6e-07 AD=2.24e-14 AS=1.84e-14 PD=6e-07 PS=5.5e-07 $X=127300 $Y=55775 $D=0
M1135 398 386 VDD VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=2.24e-14 AS=1.84e-14 PD=6e-07 PS=5.5e-07 $X=127300 $Y=58855 $D=0
M1136 205 389 396 205 PMOS_VTL L=5e-08 W=1.6e-07 AD=2.24e-14 AS=2.24e-14 PD=6e-07 PS=6e-07 $X=127680 $Y=55775 $D=0
M1137 VDD 389 398 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=2.24e-14 AS=2.24e-14 PD=6e-07 PS=6e-07 $X=127680 $Y=58855 $D=0
M1138 407 RESET 194 407 PMOS_VTL L=5e-08 W=1.6e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 $X=127905 $Y=50125 $D=0
M1139 396 166 205 205 PMOS_VTL L=5e-08 W=1.6e-07 AD=1.84e-14 AS=2.24e-14 PD=5.5e-07 PS=6e-07 $X=128060 $Y=55775 $D=0
M1140 398 167 VDD VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=1.84e-14 AS=2.24e-14 PD=5.5e-07 PS=6e-07 $X=128060 $Y=58855 $D=0
M1141 407 192 193 407 PMOS_VTL L=5e-08 W=1.6e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 $X=128765 $Y=50125 $D=0
M1142 399 195 396 205 PMOS_VTL L=5e-08 W=1.4e-07 AD=1.68e-14 AS=1.75e-14 PD=5.2e-07 PS=5.3e-07 $X=128800 $Y=55775 $D=0
M1143 400 196 398 VDD PMOS_VTL L=5e-08 W=1.4e-07 AD=1.68e-14 AS=1.75e-14 PD=5.2e-07 PS=5.3e-07 $X=128800 $Y=58855 $D=0
M1144 494 166 399 205 PMOS_VTL L=5e-08 W=1.6e-07 AD=2.24e-14 AS=1.84e-14 PD=6e-07 PS=5.5e-07 $X=129530 $Y=55775 $D=0
M1145 495 167 400 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=2.24e-14 AS=1.84e-14 PD=6e-07 PS=5.5e-07 $X=129530 $Y=58855 $D=0
M1146 407 18 192 407 PMOS_VTL L=5e-08 W=1.6e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 $X=129625 $Y=50125 $D=0
M1147 496 386 494 205 PMOS_VTL L=5e-08 W=1.6e-07 AD=2.24e-14 AS=2.24e-14 PD=6e-07 PS=6e-07 $X=129910 $Y=55775 $D=0
M1148 497 386 495 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=2.24e-14 AS=2.24e-14 PD=6e-07 PS=6e-07 $X=129910 $Y=58855 $D=0
M1149 205 389 496 205 PMOS_VTL L=5e-08 W=1.6e-07 AD=1.84e-14 AS=2.24e-14 PD=5.5e-07 PS=6e-07 $X=130290 $Y=55775 $D=0
M1150 VDD 389 497 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=1.84e-14 AS=2.24e-14 PD=5.5e-07 PS=6e-07 $X=130290 $Y=58855 $D=0
M1151 204 192 183 407 PMOS_VTL L=5e-08 W=1.6e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 $X=130485 $Y=50125 $D=0
M1152 VDD 202 389 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 $X=130920 $Y=62980 $D=0
M1153 VDD 202 201 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 $X=130920 $Y=63840 $D=0
M1154 202 201 206 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=2.4e-14 AS=1.92e-14 PD=6.2e-07 PS=5.6e-07 $X=130920 $Y=64700 $D=0
M1155 206 199 202 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=2.4e-14 AS=2.4e-14 PD=6.2e-07 PS=6.2e-07 $X=130920 $Y=65100 $D=0
M1156 VDD 197 206 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=1.92e-14 AS=2.4e-14 PD=5.6e-07 PS=6.2e-07 $X=130920 $Y=65500 $D=0
M1157 VDD RESET 199 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 $X=130920 $Y=66360 $D=0
M1158 VDD 198 197 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 $X=130920 $Y=67220 $D=0
M1159 VDD 18 198 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 $X=130920 $Y=68080 $D=0
M1160 203 198 202 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 $X=130920 $Y=68940 $D=0
M1161 498 198 VDD VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=2.24e-14 AS=1.92e-14 PD=6e-07 PS=5.6e-07 $X=130920 $Y=69800 $D=0
M1162 200 203 498 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=1.92e-14 AS=2.24e-14 PD=5.6e-07 PS=6e-07 $X=130920 $Y=70180 $D=0
M1163 203 199 VDD VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=2.4e-14 AS=1.92e-14 PD=6.2e-07 PS=5.6e-07 $X=130920 $Y=71040 $D=0
M1164 VDD 200 203 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=1.92e-14 AS=2.4e-14 PD=5.6e-07 PS=6.2e-07 $X=130920 $Y=71440 $D=0
M1165 401 197 200 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 $X=130920 $Y=72300 $D=0
M1166 VDD 402 401 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 $X=130920 $Y=73160 $D=0
M1167 VDD B6 402 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 $X=130920 $Y=74020 $D=0
M1168 499 192 407 407 PMOS_VTL L=5e-08 W=1.6e-07 AD=2.24e-14 AS=1.92e-14 PD=6e-07 PS=5.6e-07 $X=131345 $Y=50125 $D=0
M1169 VDD 400 208 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 $X=131390 $Y=58455 $D=0
M1170 404 121 205 205 PMOS_VTL L=5e-08 W=1.6e-07 AD=1.84e-14 AS=1.84e-14 PD=5.5e-07 PS=5.5e-07 $X=131420 $Y=56315 $D=0
M1171 207 204 499 407 PMOS_VTL L=5e-08 W=1.6e-07 AD=1.92e-14 AS=2.24e-14 PD=5.6e-07 PS=6e-07 $X=131725 $Y=50125 $D=0
M1172 209 121 208 205 PMOS_VTL L=5e-08 W=1.6e-07 AD=2.24e-14 AS=1.84e-14 PD=6e-07 PS=5.5e-07 $X=132190 $Y=56315 $D=0
M1173 210 399 205 205 PMOS_VTL L=5e-08 W=1.6e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 $X=132285 $Y=55135 $D=0
M1174 210 404 209 205 PMOS_VTL L=5e-08 W=1.6e-07 AD=1.84e-14 AS=2.24e-14 PD=5.5e-07 PS=6e-07 $X=132570 $Y=56315 $D=0
M1175 204 194 407 407 PMOS_VTL L=5e-08 W=1.6e-07 AD=2.4e-14 AS=1.92e-14 PD=6.2e-07 PS=5.6e-07 $X=132585 $Y=50125 $D=0
M1176 407 207 204 407 PMOS_VTL L=5e-08 W=1.6e-07 AD=1.92e-14 AS=2.4e-14 PD=5.6e-07 PS=6.2e-07 $X=132985 $Y=50125 $D=0
M1177 405 193 207 407 PMOS_VTL L=5e-08 W=1.6e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 $X=133845 $Y=50125 $D=0
M1178 407 406 405 407 PMOS_VTL L=5e-08 W=1.6e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 $X=134705 $Y=50125 $D=0
M1179 407 209 406 407 PMOS_VTL L=5e-08 W=1.6e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 $X=135565 $Y=50125 $D=0
M1180 427 409 415 427 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=2.07e-14 PD=6.4e-07 PS=5.9e-07 $X=136860 $Y=55775 $D=0
M1181 VDD 409 417 VDD PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=2.07e-14 PD=6.4e-07 PS=5.9e-07 $X=136860 $Y=58855 $D=0
M1182 433 218 S7 433 PMOS_VTL L=5e-08 W=1.6e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 $X=136905 $Y=50125 $D=0
M1183 VDD 410 409 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 $X=137115 $Y=61795 $D=0
M1184 VDD 216 410 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 $X=137125 $Y=62980 $D=0
M1185 VDD 216 215 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 $X=137125 $Y=63840 $D=0
M1186 216 215 219 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=2.4e-14 AS=1.92e-14 PD=6.2e-07 PS=5.6e-07 $X=137125 $Y=64700 $D=0
M1187 219 213 216 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=2.4e-14 AS=2.4e-14 PD=6.2e-07 PS=6.2e-07 $X=137125 $Y=65100 $D=0
M1188 VDD 211 219 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=1.92e-14 AS=2.4e-14 PD=5.6e-07 PS=6.2e-07 $X=137125 $Y=65500 $D=0
M1189 VDD RESET 213 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 $X=137125 $Y=66360 $D=0
M1190 VDD 212 211 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 $X=137125 $Y=67220 $D=0
M1191 VDD 18 212 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 $X=137125 $Y=68080 $D=0
M1192 217 212 216 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 $X=137125 $Y=68940 $D=0
M1193 500 212 VDD VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=2.24e-14 AS=1.92e-14 PD=6e-07 PS=5.6e-07 $X=137125 $Y=69800 $D=0
M1194 214 217 500 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=1.92e-14 AS=2.24e-14 PD=5.6e-07 PS=6e-07 $X=137125 $Y=70180 $D=0
M1195 217 213 VDD VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=2.4e-14 AS=1.92e-14 PD=6.2e-07 PS=5.6e-07 $X=137125 $Y=71040 $D=0
M1196 VDD 214 217 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=1.92e-14 AS=2.4e-14 PD=5.6e-07 PS=6.2e-07 $X=137125 $Y=71440 $D=0
M1197 411 211 214 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 $X=137125 $Y=72300 $D=0
M1198 VDD 412 411 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 $X=137125 $Y=73160 $D=0
M1199 VDD A7 412 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 $X=137125 $Y=74020 $D=0
M1200 415 413 427 427 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=2.52e-14 PD=6.4e-07 PS=6.4e-07 $X=137240 $Y=55775 $D=0
M1201 417 413 VDD VDD PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=2.52e-14 PD=6.4e-07 PS=6.4e-07 $X=137240 $Y=58855 $D=0
M1202 225 195 415 427 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=2.52e-14 PD=6.4e-07 PS=6.4e-07 $X=137620 $Y=55775 $D=0
M1203 226 196 417 VDD PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=2.52e-14 PD=6.4e-07 PS=6.4e-07 $X=137620 $Y=58855 $D=0
M1204 433 218 220 433 PMOS_VTL L=5e-08 W=1.6e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 $X=137765 $Y=50125 $D=0
M1205 501 409 225 427 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=2.52e-14 PD=6.4e-07 PS=6.4e-07 $X=138000 $Y=55775 $D=0
M1206 502 409 226 VDD PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=2.52e-14 PD=6.4e-07 PS=6.4e-07 $X=138000 $Y=58855 $D=0
M1207 427 413 501 427 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.07e-14 AS=2.52e-14 PD=5.9e-07 PS=6.4e-07 $X=138380 $Y=55775 $D=0
M1208 VDD 413 502 VDD PMOS_VTL L=5e-08 W=1.8e-07 AD=2.07e-14 AS=2.52e-14 PD=5.9e-07 PS=6.4e-07 $X=138380 $Y=58855 $D=0
M1209 218 220 221 433 PMOS_VTL L=5e-08 W=1.6e-07 AD=2.4e-14 AS=1.92e-14 PD=6.2e-07 PS=5.6e-07 $X=138625 $Y=50125 $D=0
M1210 221 224 218 433 PMOS_VTL L=5e-08 W=1.6e-07 AD=2.4e-14 AS=2.4e-14 PD=6.2e-07 PS=6.2e-07 $X=139025 $Y=50125 $D=0
M1211 420 409 427 427 PMOS_VTL L=5e-08 W=1.6e-07 AD=2.24e-14 AS=1.84e-14 PD=6e-07 PS=5.5e-07 $X=139100 $Y=55775 $D=0
M1212 422 409 VDD VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=2.24e-14 AS=1.84e-14 PD=6e-07 PS=5.5e-07 $X=139100 $Y=58855 $D=0
M1213 433 223 221 433 PMOS_VTL L=5e-08 W=1.6e-07 AD=1.92e-14 AS=2.4e-14 PD=5.6e-07 PS=6.2e-07 $X=139425 $Y=50125 $D=0
M1214 427 413 420 427 PMOS_VTL L=5e-08 W=1.6e-07 AD=2.24e-14 AS=2.24e-14 PD=6e-07 PS=6e-07 $X=139480 $Y=55775 $D=0
M1215 VDD 413 422 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=2.24e-14 AS=2.24e-14 PD=6e-07 PS=6e-07 $X=139480 $Y=58855 $D=0
M1216 420 195 427 427 PMOS_VTL L=5e-08 W=1.6e-07 AD=1.84e-14 AS=2.24e-14 PD=5.5e-07 PS=6e-07 $X=139860 $Y=55775 $D=0
M1217 422 196 VDD VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=1.84e-14 AS=2.24e-14 PD=5.5e-07 PS=6e-07 $X=139860 $Y=58855 $D=0
M1218 433 RESET 224 433 PMOS_VTL L=5e-08 W=1.6e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 $X=140285 $Y=50125 $D=0
M1219 423 225 420 427 PMOS_VTL L=5e-08 W=1.4e-07 AD=1.68e-14 AS=1.75e-14 PD=5.2e-07 PS=5.3e-07 $X=140600 $Y=55775 $D=0
M1220 236 226 422 VDD PMOS_VTL L=5e-08 W=1.4e-07 AD=1.68e-14 AS=1.75e-14 PD=5.2e-07 PS=5.3e-07 $X=140600 $Y=58855 $D=0
M1221 433 222 223 433 PMOS_VTL L=5e-08 W=1.6e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 $X=141145 $Y=50125 $D=0
M1222 503 195 423 427 PMOS_VTL L=5e-08 W=1.6e-07 AD=2.24e-14 AS=1.84e-14 PD=6e-07 PS=5.5e-07 $X=141330 $Y=55775 $D=0
M1223 504 196 236 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=2.24e-14 AS=1.84e-14 PD=6e-07 PS=5.5e-07 $X=141330 $Y=58855 $D=0
M1224 505 409 503 427 PMOS_VTL L=5e-08 W=1.6e-07 AD=2.24e-14 AS=2.24e-14 PD=6e-07 PS=6e-07 $X=141710 $Y=55775 $D=0
M1225 506 409 504 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=2.24e-14 AS=2.24e-14 PD=6e-07 PS=6e-07 $X=141710 $Y=58855 $D=0
M1226 433 18 222 433 PMOS_VTL L=5e-08 W=1.6e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 $X=142005 $Y=50125 $D=0
M1227 427 413 505 427 PMOS_VTL L=5e-08 W=1.6e-07 AD=1.84e-14 AS=2.24e-14 PD=5.5e-07 PS=6e-07 $X=142090 $Y=55775 $D=0
M1228 VDD 413 506 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=1.84e-14 AS=2.24e-14 PD=5.5e-07 PS=6e-07 $X=142090 $Y=58855 $D=0
M1229 VDD 424 413 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 $X=142635 $Y=61795 $D=0
M1230 VDD 232 424 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 $X=142645 $Y=62980 $D=0
M1231 VDD 232 231 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 $X=142645 $Y=63840 $D=0
M1232 232 231 234 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=2.4e-14 AS=1.92e-14 PD=6.2e-07 PS=5.6e-07 $X=142645 $Y=64700 $D=0
M1233 234 229 232 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=2.4e-14 AS=2.4e-14 PD=6.2e-07 PS=6.2e-07 $X=142645 $Y=65100 $D=0
M1234 VDD 227 234 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=1.92e-14 AS=2.4e-14 PD=5.6e-07 PS=6.2e-07 $X=142645 $Y=65500 $D=0
M1235 VDD RESET 229 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 $X=142645 $Y=66360 $D=0
M1236 VDD 228 227 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 $X=142645 $Y=67220 $D=0
M1237 VDD 18 228 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 $X=142645 $Y=68080 $D=0
M1238 233 228 232 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 $X=142645 $Y=68940 $D=0
M1239 507 228 VDD VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=2.24e-14 AS=1.92e-14 PD=6e-07 PS=5.6e-07 $X=142645 $Y=69800 $D=0
M1240 230 233 507 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=1.92e-14 AS=2.24e-14 PD=5.6e-07 PS=6e-07 $X=142645 $Y=70180 $D=0
M1241 233 229 VDD VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=2.4e-14 AS=1.92e-14 PD=6.2e-07 PS=5.6e-07 $X=142645 $Y=71040 $D=0
M1242 VDD 230 233 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=1.92e-14 AS=2.4e-14 PD=5.6e-07 PS=6.2e-07 $X=142645 $Y=71440 $D=0
M1243 425 227 230 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 $X=142645 $Y=72300 $D=0
M1244 VDD 426 425 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 $X=142645 $Y=73160 $D=0
M1245 VDD B7 426 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 $X=142645 $Y=74020 $D=0
M1246 235 222 218 433 PMOS_VTL L=5e-08 W=1.6e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 $X=142865 $Y=50125 $D=0
M1247 429 121 427 427 PMOS_VTL L=5e-08 W=1.6e-07 AD=1.84e-14 AS=1.84e-14 PD=5.5e-07 PS=5.5e-07 $X=143220 $Y=56315 $D=0
M1248 508 222 433 433 PMOS_VTL L=5e-08 W=1.6e-07 AD=2.24e-14 AS=1.92e-14 PD=6e-07 PS=5.6e-07 $X=143725 $Y=50125 $D=0
M1249 237 121 236 427 PMOS_VTL L=5e-08 W=1.6e-07 AD=2.24e-14 AS=1.84e-14 PD=6e-07 PS=5.5e-07 $X=143990 $Y=56315 $D=0
M1250 238 235 508 433 PMOS_VTL L=5e-08 W=1.6e-07 AD=1.92e-14 AS=2.24e-14 PD=5.6e-07 PS=6e-07 $X=144105 $Y=50125 $D=0
M1251 239 429 237 427 PMOS_VTL L=5e-08 W=1.6e-07 AD=1.84e-14 AS=2.24e-14 PD=5.5e-07 PS=6e-07 $X=144370 $Y=56315 $D=0
M1252 235 224 433 433 PMOS_VTL L=5e-08 W=1.6e-07 AD=2.4e-14 AS=1.92e-14 PD=6.2e-07 PS=5.6e-07 $X=144965 $Y=50125 $D=0
M1253 433 238 235 433 PMOS_VTL L=5e-08 W=1.6e-07 AD=1.92e-14 AS=2.4e-14 PD=5.6e-07 PS=6.2e-07 $X=145365 $Y=50125 $D=0
M1254 431 223 238 433 PMOS_VTL L=5e-08 W=1.6e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 $X=146225 $Y=50125 $D=0
M1255 430 121 VDD VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=1.84e-14 AS=1.84e-14 PD=5.5e-07 PS=5.5e-07 $X=146325 $Y=56290 $D=0
M1256 433 432 431 433 PMOS_VTL L=5e-08 W=1.6e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 $X=147085 $Y=50125 $D=0
M1257 VDD 121 226 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=2.24e-14 AS=1.84e-14 PD=6e-07 PS=5.5e-07 $X=147095 $Y=56290 $D=0
M1258 225 430 VDD VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=1.84e-14 AS=2.24e-14 PD=5.5e-07 PS=6e-07 $X=147475 $Y=56290 $D=0
M1259 433 237 432 433 PMOS_VTL L=5e-08 W=1.6e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 $X=147945 $Y=50125 $D=0
M1260 435 VDD VDD VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 $X=149095 $Y=57685 $D=0
M1261 436 435 VDD VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 $X=149095 $Y=58545 $D=0
M1262 246 240 436 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 $X=149095 $Y=59405 $D=0
M1263 247 246 VDD VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=2.4e-14 AS=1.92e-14 PD=6.2e-07 PS=5.6e-07 $X=149095 $Y=60265 $D=0
M1264 VDD 243 247 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=1.92e-14 AS=2.4e-14 PD=5.6e-07 PS=6.2e-07 $X=149095 $Y=60665 $D=0
M1265 509 247 246 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=2.24e-14 AS=1.92e-14 PD=6e-07 PS=5.6e-07 $X=149095 $Y=61525 $D=0
M1266 VDD 244 509 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=1.92e-14 AS=2.24e-14 PD=5.6e-07 PS=6e-07 $X=149095 $Y=61905 $D=0
M1267 242 244 247 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 $X=149095 $Y=62765 $D=0
M1268 244 18 VDD VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 $X=149095 $Y=63625 $D=0
M1269 240 244 VDD VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 $X=149095 $Y=64485 $D=0
M1270 243 RESET VDD VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 $X=149095 $Y=65345 $D=0
M1271 245 240 VDD VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=2.4e-14 AS=1.92e-14 PD=6.2e-07 PS=5.6e-07 $X=149095 $Y=66205 $D=0
M1272 242 243 245 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=2.4e-14 AS=2.4e-14 PD=6.2e-07 PS=6.2e-07 $X=149095 $Y=66605 $D=0
M1273 245 241 242 VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=1.92e-14 AS=2.4e-14 PD=5.6e-07 PS=6.2e-07 $X=149095 $Y=67005 $D=0
M1274 241 242 VDD VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 $X=149095 $Y=67865 $D=0
M1275 434 242 VDD VDD PMOS_VTL L=5e-08 W=1.6e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 $X=149095 $Y=68725 $D=0
.ENDS
***************************************
